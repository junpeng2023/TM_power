module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in3,
    in4,
    in5,
    in6,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out3,
    out4,
    out5,
    out6,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in3;
 input in4;
 input in5;
 input in6;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out3;
 output out4;
 output out5;
 output out6;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net363;
 wire net785;
 wire net800;
 wire net833;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net931;
 wire clknet_1_0__leaf_net931;
 wire clknet_1_1__leaf_net931;
 wire clknet_0_net329;
 wire clknet_1_0__leaf_net329;
 wire clknet_1_1__leaf_net329;
 wire clknet_0_net985;
 wire clknet_1_0__leaf_net985;
 wire clknet_1_1__leaf_net985;
 wire clknet_0_net361;
 wire clknet_1_0__leaf_net361;
 wire clknet_1_1__leaf_net361;
 wire clknet_0_net830;
 wire clknet_1_0__leaf_net830;
 wire clknet_1_1__leaf_net830;
 wire clknet_0_net338;
 wire clknet_1_0__leaf_net338;
 wire clknet_1_1__leaf_net338;
 wire clknet_0_net983;
 wire clknet_1_0__leaf_net983;
 wire clknet_1_1__leaf_net983;
 wire clknet_0_net292;
 wire clknet_1_0__leaf_net292;
 wire clknet_1_1__leaf_net292;
 wire clknet_0_net427;
 wire clknet_1_0__leaf_net427;
 wire clknet_1_1__leaf_net427;
 wire clknet_0_net929;
 wire clknet_1_0__leaf_net929;
 wire clknet_1_1__leaf_net929;
 wire clknet_0_net447;
 wire clknet_1_0__leaf_net447;
 wire clknet_1_1__leaf_net447;
 wire clknet_0_net930;
 wire clknet_1_0__leaf_net930;
 wire clknet_1_1__leaf_net930;
 wire clknet_0_net451;
 wire clknet_1_0__leaf_net451;
 wire clknet_1_1__leaf_net451;
 wire clknet_0_net481;
 wire clknet_1_0__leaf_net481;
 wire clknet_1_1__leaf_net481;
 wire clknet_0_net719;
 wire clknet_1_0__leaf_net719;
 wire clknet_1_1__leaf_net719;
 wire clknet_0_net593;
 wire clknet_1_0__leaf_net593;
 wire clknet_1_1__leaf_net593;
 wire clknet_0_net458;
 wire clknet_1_0__leaf_net458;
 wire clknet_1_1__leaf_net458;
 wire clknet_0_net448;
 wire clknet_1_0__leaf_net448;
 wire clknet_1_1__leaf_net448;
 wire clknet_0_net877;
 wire clknet_1_0__leaf_net877;
 wire clknet_1_1__leaf_net877;
 wire clknet_0_net894;
 wire clknet_1_0__leaf_net894;
 wire clknet_1_1__leaf_net894;
 wire clknet_0_net605;
 wire clknet_1_0__leaf_net605;
 wire clknet_1_1__leaf_net605;
 wire clknet_0_net567;
 wire clknet_1_0__leaf_net567;
 wire clknet_1_1__leaf_net567;
 wire clknet_0_net609;
 wire clknet_1_0__leaf_net609;
 wire clknet_1_1__leaf_net609;
 wire clknet_0_net449;
 wire clknet_1_0__leaf_net449;
 wire clknet_1_1__leaf_net449;
 wire clknet_0_net457;
 wire clknet_1_0__leaf_net457;
 wire clknet_1_1__leaf_net457;
 wire clknet_0_net911;
 wire clknet_1_0__leaf_net911;
 wire clknet_1_1__leaf_net911;
 wire clknet_0_net707;
 wire clknet_1_0__leaf_net707;
 wire clknet_1_1__leaf_net707;
 wire clknet_0_net452;
 wire clknet_1_0__leaf_net452;
 wire clknet_1_1__leaf_net452;
 wire clknet_0_net463;
 wire clknet_1_0__leaf_net463;
 wire clknet_1_1__leaf_net463;
 wire clknet_0_net821;
 wire clknet_1_0__leaf_net821;
 wire clknet_1_1__leaf_net821;
 wire clknet_0_net546;
 wire clknet_1_0__leaf_net546;
 wire clknet_1_1__leaf_net546;
 wire clknet_0_net876;
 wire clknet_1_0__leaf_net876;
 wire clknet_1_1__leaf_net876;
 wire clknet_0_net436;
 wire clknet_1_0__leaf_net436;
 wire clknet_1_1__leaf_net436;
 wire clknet_0_net895;
 wire clknet_1_0__leaf_net895;
 wire clknet_1_1__leaf_net895;
 wire clknet_0_net913;
 wire clknet_1_0__leaf_net913;
 wire clknet_1_1__leaf_net913;
 wire clknet_0_net709;
 wire clknet_1_0__leaf_net709;
 wire clknet_1_1__leaf_net709;
 wire clknet_0_net912;
 wire clknet_1_0__leaf_net912;
 wire clknet_1_1__leaf_net912;
 wire clknet_0_net893;
 wire clknet_1_0__leaf_net893;
 wire clknet_1_1__leaf_net893;
 wire clknet_0_net875;
 wire clknet_1_0__leaf_net875;
 wire clknet_1_1__leaf_net875;
 wire clknet_0_net420;
 wire clknet_1_0__leaf_net420;
 wire clknet_1_1__leaf_net420;
 wire clknet_0_net464;
 wire clknet_1_0__leaf_net464;
 wire clknet_1_1__leaf_net464;
 wire clknet_0_net424;
 wire clknet_1_0__leaf_net424;
 wire clknet_1_1__leaf_net424;
 wire clknet_0_net856;
 wire clknet_1_0__leaf_net856;
 wire clknet_1_1__leaf_net856;
 wire clknet_0_net353;
 wire clknet_1_0__leaf_net353;
 wire clknet_1_1__leaf_net353;
 wire clknet_0_net221;
 wire clknet_1_0__leaf_net221;
 wire clknet_1_1__leaf_net221;
 wire clknet_0_net855;
 wire clknet_1_0__leaf_net855;
 wire clknet_1_1__leaf_net855;
 wire clknet_0_net823;
 wire clknet_1_0__leaf_net823;
 wire clknet_1_1__leaf_net823;
 wire clknet_0_net346;
 wire clknet_1_0__leaf_net346;
 wire clknet_1_1__leaf_net346;
 wire clknet_0_net974;
 wire clknet_1_0__leaf_net974;
 wire clknet_1_1__leaf_net974;
 wire clknet_0_net354;
 wire clknet_1_0__leaf_net354;
 wire clknet_1_1__leaf_net354;
 wire clknet_0_net854;
 wire clknet_1_0__leaf_net854;
 wire clknet_1_1__leaf_net854;
 wire clknet_0_net969;
 wire clknet_1_0__leaf_net969;
 wire clknet_1_1__leaf_net969;
 wire clknet_0_net315;
 wire clknet_1_0__leaf_net315;
 wire clknet_1_1__leaf_net315;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;

 sky130_fd_sc_hd__and2_1 c100 (.A(net68),
    .B(net850),
    .X(net74));
 sky130_fd_sc_hd__and2_1 c101 (.A(net50),
    .B(net851),
    .X(net75));
 sky130_fd_sc_hd__and2_0 c102 (.A(net75),
    .B(net67),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 c103 (.A(net802),
    .X(net77));
 sky130_fd_sc_hd__dlymetal6s2s_1 c104 (.A(net766),
    .X(net78));
 sky130_fd_sc_hd__dlymetal6s2s_1 c105 (.A(net802),
    .X(net973));
 sky130_fd_sc_hd__and3_2 c106 (.A(net67),
    .B(net973),
    .C(net1051),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 c107 (.A(net802),
    .X(net80));
 sky130_fd_sc_hd__and3_2 c108 (.A(net77),
    .B(net73),
    .C(net80),
    .X(net81));
 sky130_fd_sc_hd__mux4_1 c109 (.A0(net80),
    .A1(net76),
    .A2(net79),
    .A3(net81),
    .S0(net1011),
    .S1(net847),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 c110 (.A(net819),
    .X(net83));
 sky130_fd_sc_hd__and2_1 c111 (.A(net6),
    .B(net81),
    .X(net84));
 sky130_fd_sc_hd__dlymetal6s2s_1 c112 (.A(net818),
    .X(net85));
 sky130_fd_sc_hd__and2_1 c113 (.A(net37),
    .B(net851),
    .X(net86));
 sky130_fd_sc_hd__and2_1 c114 (.A(net946),
    .B(net85),
    .X(net87));
 sky130_fd_sc_hd__and2_1 c115 (.A(net973),
    .B(net962),
    .X(net88));
 sky130_fd_sc_hd__and3_1 c116 (.A(net35),
    .B(net37),
    .C(net86),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 c117 (.A(net756),
    .X(net90));
 sky130_fd_sc_hd__and2_0 c118 (.A(net86),
    .B(net848),
    .X(net91));
 sky130_fd_sc_hd__and2_1 c119 (.A(net87),
    .B(net85),
    .X(net92));
 sky130_fd_sc_hd__and2_2 c120 (.A(net85),
    .B(net92),
    .X(net93));
 sky130_fd_sc_hd__and2_0 c121 (.A(net31),
    .B(net92),
    .X(net94));
 sky130_fd_sc_hd__and3_1 c122 (.A(net90),
    .B(net86),
    .C(net84),
    .X(net95));
 sky130_fd_sc_hd__and2_2 c123 (.A(net86),
    .B(net85),
    .X(net96));
 sky130_fd_sc_hd__and2_0 c124 (.A(net92),
    .B(net87),
    .X(net97));
 sky130_fd_sc_hd__mux4_1 c125 (.A0(net23),
    .A1(net85),
    .A2(net96),
    .A3(net15),
    .S0(net79),
    .S1(net68),
    .X(net98));
 sky130_fd_sc_hd__buf_2 c126 (.A(net766),
    .X(net99));
 sky130_fd_sc_hd__mux4_1 c127 (.A0(net83),
    .A1(net87),
    .A2(net92),
    .A3(net96),
    .S0(net85),
    .S1(net75),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 c128 (.A(net802),
    .X(net101));
 sky130_fd_sc_hd__and2_0 c129 (.A(net94),
    .B(net81),
    .X(net102));
 sky130_fd_sc_hd__or4bb_1 c130 (.A(net102),
    .B(net99),
    .C_N(net85),
    .D_N(net88),
    .X(net103));
 sky130_fd_sc_hd__mux4_1 c131 (.A0(net103),
    .A1(net92),
    .A2(net86),
    .A3(net68),
    .S0(net851),
    .S1(net1007),
    .X(net104));
 sky130_fd_sc_hd__and2_1 c132 (.A(net963),
    .B(net955),
    .X(net105));
 sky130_fd_sc_hd__and2_2 c133 (.A(net363),
    .B(net947),
    .X(net106));
 sky130_fd_sc_hd__and2_4 c134 (.A(net946),
    .B(net955),
    .X(net107));
 sky130_fd_sc_hd__and2_2 c135 (.A(net949),
    .B(net107),
    .X(net108));
 sky130_fd_sc_hd__and3_2 c136 (.A(net800),
    .B(net947),
    .C(net963),
    .X(net109));
 sky130_fd_sc_hd__and2_1 c137 (.A(net109),
    .B(net107),
    .X(net110));
 sky130_fd_sc_hd__and2_2 c138 (.A(net108),
    .B(net785),
    .X(net111));
 sky130_fd_sc_hd__and2_2 c139 (.A(net959),
    .B(net833),
    .X(net112));
 sky130_fd_sc_hd__and2_1 c140 (.A(net947),
    .B(net107),
    .X(net113));
 sky130_fd_sc_hd__and2_4 c141 (.A(net112),
    .B(net111),
    .X(net114));
 sky130_fd_sc_hd__or4bb_4 c142 (.A(net111),
    .B(net105),
    .C_N(net113),
    .D_N(net114),
    .X(net115));
 sky130_fd_sc_hd__and3_1 c143 (.A(net959),
    .B(net113),
    .C(net114),
    .X(net116));
 sky130_fd_sc_hd__or4bb_4 c144 (.A(net109),
    .B(net115),
    .C_N(net116),
    .D_N(net111),
    .X(net117));
 sky130_fd_sc_hd__and2_2 c145 (.A(net785),
    .B(net116),
    .X(net118));
 sky130_fd_sc_hd__a2111o_4 c146 (.A1(net116),
    .A2(net118),
    .B1(net110),
    .C1(net108),
    .D1(net109),
    .X(net119));
 sky130_fd_sc_hd__a2111o_2 c147 (.A1(net116),
    .A2(net111),
    .B1(net115),
    .C1(net109),
    .D1(net959),
    .X(net120));
 sky130_fd_sc_hd__a2111o_4 c148 (.A1(net115),
    .A2(net119),
    .B1(net109),
    .C1(net110),
    .D1(net120),
    .X(net986));
 sky130_fd_sc_hd__and3_2 c149 (.A(net105),
    .B(net107),
    .C(net118),
    .X(net121));
 sky130_fd_sc_hd__and2_2 c150 (.A(net121),
    .B(net949),
    .X(net122));
 sky130_fd_sc_hd__and3_1 c151 (.A(net117),
    .B(net121),
    .C(net122),
    .X(net123));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net122),
    .A1(net123),
    .A2(net120),
    .A3(net121),
    .S0(net107),
    .S1(net115),
    .X(net124));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net123),
    .A1(net106),
    .A2(net959),
    .A3(net105),
    .S0(net124),
    .S1(net122),
    .X(net125));
 sky130_fd_sc_hd__and2_2 c154 (.A(net946),
    .B(net950),
    .X(net126));
 sky130_fd_sc_hd__and3_2 c155 (.A(net833),
    .B(net126),
    .C(net2),
    .X(net127));
 sky130_fd_sc_hd__and2_1 c156 (.A(net800),
    .B(net2),
    .X(net128));
 sky130_fd_sc_hd__and2_1 c157 (.A(net948),
    .B(net958),
    .X(net129));
 sky130_fd_sc_hd__or4bb_4 c158 (.A(net127),
    .B(net108),
    .C_N(net126),
    .D_N(net119),
    .X(net130));
 sky130_fd_sc_hd__and2_2 c159 (.A(net3),
    .B(net130),
    .X(net131));
 sky130_fd_sc_hd__and2_1 c160 (.A(net952),
    .B(net956),
    .X(net132));
 sky130_fd_sc_hd__or4bb_1 c161 (.A(net961),
    .B(net5),
    .C_N(net107),
    .D_N(net115),
    .X(net133));
 sky130_fd_sc_hd__and2_1 c162 (.A(net128),
    .B(net130),
    .X(net134));
 sky130_fd_sc_hd__and2_4 c163 (.A(net16),
    .B(net132),
    .X(net135));
 sky130_fd_sc_hd__mux4_2 c164 (.A0(net133),
    .A1(net945),
    .A2(net135),
    .A3(net134),
    .S0(net958),
    .S1(net128),
    .X(net136));
 sky130_fd_sc_hd__or4bb_2 c165 (.A(net133),
    .B(net961),
    .C_N(net950),
    .D_N(net953),
    .X(net137));
 sky130_fd_sc_hd__a2111o_1 c166 (.A1(net958),
    .A2(net117),
    .B1(net132),
    .C1(net114),
    .D1(net129),
    .X(net138));
 sky130_fd_sc_hd__or4bb_4 c167 (.A(net17),
    .B(net129),
    .C_N(net138),
    .D_N(net946),
    .X(net139));
 sky130_fd_sc_hd__and3_1 c168 (.A(net6),
    .B(net16),
    .C(net127),
    .X(net140));
 sky130_fd_sc_hd__and2_1 c169 (.A(net8),
    .B(net134),
    .X(net141));
 sky130_fd_sc_hd__a2111o_4 c170 (.A1(net135),
    .A2(net16),
    .B1(net5),
    .C1(net137),
    .D1(net139),
    .X(net142));
 sky130_fd_sc_hd__or4bb_1 c171 (.A(net139),
    .B(net132),
    .C_N(net133),
    .D_N(net1001),
    .X(net143));
 sky130_fd_sc_hd__or4bb_2 c172 (.A(net136),
    .B(net129),
    .C_N(net956),
    .D_N(net1001),
    .X(net144));
 sky130_fd_sc_hd__a2111o_4 c173 (.A1(net141),
    .A2(net127),
    .B1(net138),
    .C1(net958),
    .D1(net1001),
    .X(net145));
 sky130_fd_sc_hd__and3_1 c174 (.A(net136),
    .B(net140),
    .C(net137),
    .X(net146));
 sky130_fd_sc_hd__and2_2 c175 (.A(net146),
    .B(net363),
    .X(net147));
 sky130_fd_sc_hd__and2_1 c176 (.A(net27),
    .B(net131),
    .X(net148));
 sky130_fd_sc_hd__and2_1 c177 (.A(net148),
    .B(net143),
    .X(net149));
 sky130_fd_sc_hd__and2_1 c178 (.A(net14),
    .B(net135),
    .X(net150));
 sky130_fd_sc_hd__and2_1 c179 (.A(net998),
    .B(net108),
    .X(net151));
 sky130_fd_sc_hd__and2_0 c180 (.A(net1032),
    .B(net148),
    .X(net152));
 sky130_fd_sc_hd__and3_1 c181 (.A(net152),
    .B(net148),
    .C(net8),
    .X(net153));
 sky130_fd_sc_hd__and3_1 c182 (.A(net33),
    .B(net27),
    .C(net1031),
    .X(net154));
 sky130_fd_sc_hd__and2_1 c183 (.A(net30),
    .B(net21),
    .X(net155));
 sky130_fd_sc_hd__and2_4 c184 (.A(net135),
    .B(net33),
    .X(net156));
 sky130_fd_sc_hd__and2_2 c185 (.A(net833),
    .B(net986),
    .X(net157));
 sky130_fd_sc_hd__and2_1 c186 (.A(net156),
    .B(net37),
    .X(net158));
 sky130_fd_sc_hd__mux4_2 c187 (.A0(net114),
    .A1(net156),
    .A2(net157),
    .A3(net18),
    .S0(net112),
    .S1(net135),
    .X(net159));
 sky130_fd_sc_hd__mux4_2 c188 (.A0(net138),
    .A1(net156),
    .A2(net137),
    .A3(net27),
    .S0(net148),
    .S1(net157),
    .X(net160));
 sky130_fd_sc_hd__a2111o_1 c189 (.A1(net950),
    .A2(net157),
    .B1(net156),
    .C1(net11),
    .D1(net160),
    .X(net161));
 sky130_fd_sc_hd__a2111o_4 c190 (.A1(net159),
    .A2(net124),
    .B1(net1012),
    .C1(net995),
    .D1(net156),
    .X(net162));
 sky130_fd_sc_hd__a2111o_1 c191 (.A1(net21),
    .A2(net160),
    .B1(net159),
    .C1(net33),
    .D1(net995),
    .X(net163));
 sky130_fd_sc_hd__and3_1 c192 (.A(net137),
    .B(net995),
    .C(net27),
    .X(net164));
 sky130_fd_sc_hd__a2111o_1 c193 (.A1(net143),
    .A2(net151),
    .B1(net27),
    .C1(net149),
    .D1(net995),
    .X(net165));
 sky130_fd_sc_hd__and3_1 c194 (.A(net165),
    .B(net155),
    .C(net159),
    .X(net166));
 sky130_fd_sc_hd__mux4_1 c195 (.A0(net131),
    .A1(net155),
    .A2(net1012),
    .A3(net165),
    .S0(net995),
    .S1(net137),
    .X(net167));
 sky130_fd_sc_hd__mux4_1 c196 (.A0(net157),
    .A1(net167),
    .A2(net159),
    .A3(net156),
    .S0(net148),
    .S1(net995),
    .X(net168));
 sky130_fd_sc_hd__mux4_1 c197 (.A0(net38),
    .A1(net117),
    .A2(net954),
    .A3(net995),
    .S0(net151),
    .S1(net155),
    .X(net169));
 sky130_fd_sc_hd__and2_0 c198 (.A(net140),
    .B(net106),
    .X(net170));
 sky130_fd_sc_hd__and2_2 c199 (.A(net170),
    .B(net53),
    .X(net171));
 sky130_fd_sc_hd__and2_4 c200 (.A(net127),
    .B(net45),
    .X(net172));
 sky130_fd_sc_hd__and3_1 c201 (.A(net126),
    .B(net172),
    .C(net165),
    .X(net173));
 sky130_fd_sc_hd__and3_4 c202 (.A(net156),
    .B(net972),
    .C(net163),
    .X(net174));
 sky130_fd_sc_hd__and2_0 c203 (.A(net134),
    .B(net14),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 c204 (.A(net790),
    .X(net176));
 sky130_fd_sc_hd__sdfrbp_1 c205 (.CLK(clknet_4_2_0_clk),
    .D(net171),
    .RESET_B(net46),
    .SCD(net1031),
    .SCE(net174),
    .Q(net178),
    .Q_N(net177));
 sky130_fd_sc_hd__and3_1 c206 (.A(net176),
    .B(net55),
    .C(net177),
    .X(net179));
 sky130_fd_sc_hd__and2_2 c207 (.A(net159),
    .B(net178),
    .X(net180));
 sky130_fd_sc_hd__and3_1 c208 (.A(net47),
    .B(net35),
    .C(net996),
    .X(net181));
 sky130_fd_sc_hd__and3_4 c209 (.A(net179),
    .B(net126),
    .C(net996),
    .X(net182));
 sky130_fd_sc_hd__and3_1 c210 (.A(net53),
    .B(net134),
    .C(net180),
    .X(net183));
 sky130_fd_sc_hd__and2_1 c211 (.A(net163),
    .B(net178),
    .X(net184));
 sky130_fd_sc_hd__a2111o_1 c212 (.A1(net181),
    .A2(net150),
    .B1(net177),
    .C1(net1016),
    .D1(net179),
    .X(net185));
 sky130_fd_sc_hd__buf_1 c213 (.A(net797),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 c214 (.A(net790),
    .X(net187));
 sky130_fd_sc_hd__or4bb_4 c215 (.A(net175),
    .B(net186),
    .C_N(net180),
    .D_N(net39),
    .X(net188));
 sky130_fd_sc_hd__a2111o_1 c216 (.A1(net39),
    .A2(net186),
    .B1(net157),
    .C1(net188),
    .D1(net791),
    .X(net189));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(net184),
    .A1(net189),
    .A2(net179),
    .A3(net174),
    .S0(net945),
    .S1(net177),
    .X(net190));
 sky130_fd_sc_hd__and3_4 c218 (.A(net186),
    .B(net180),
    .C(net188),
    .X(net191));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net178),
    .A1(net187),
    .A2(net182),
    .A3(net186),
    .S0(net171),
    .S1(net174),
    .X(net192));
 sky130_fd_sc_hd__and2_0 c220 (.A(net150),
    .B(net946),
    .X(net193));
 sky130_fd_sc_hd__and2_0 c221 (.A(net157),
    .B(net852),
    .X(net194));
 sky130_fd_sc_hd__or4bb_1 c222 (.A(net194),
    .B(net71),
    .C_N(net157),
    .D_N(net66),
    .X(net195));
 sky130_fd_sc_hd__and2_0 c223 (.A(net45),
    .B(clknet_1_0__leaf_net854),
    .X(net196));
 sky130_fd_sc_hd__sdfbbn_1 c224 (.CLK_N(clknet_4_8_0_clk),
    .D(net46),
    .RESET_B(net948),
    .SCD(net18),
    .SCE(net962),
    .SET_B(net996),
    .Q(net198),
    .Q_N(net197));
 sky130_fd_sc_hd__and2_0 c225 (.A(net196),
    .B(clknet_1_0__leaf_net855),
    .X(net199));
 sky130_fd_sc_hd__buf_1 c226 (.A(net726),
    .X(net200));
 sky130_fd_sc_hd__or4bb_4 c227 (.A(net69),
    .B(net997),
    .C_N(net829),
    .D_N(net1037),
    .X(net201));
 sky130_fd_sc_hd__and3_1 c228 (.A(net193),
    .B(net1018),
    .C(net829),
    .X(net202));
 sky130_fd_sc_hd__buf_1 c229 (.A(net726),
    .X(net203));
 sky130_fd_sc_hd__or4bb_1 c230 (.A(net149),
    .B(net78),
    .C_N(net174),
    .D_N(net1037),
    .X(net204));
 sky130_fd_sc_hd__sdfbbn_1 c231 (.CLK_N(clknet_4_8_0_clk),
    .D(net202),
    .RESET_B(net1025),
    .SCD(net66),
    .SCE(net69),
    .SET_B(net803),
    .Q(net206),
    .Q_N(net205));
 sky130_fd_sc_hd__mux4_1 c232 (.A0(net992),
    .A1(net203),
    .A2(net198),
    .A3(net963),
    .S0(net172),
    .S1(net803),
    .X(net207));
 sky130_fd_sc_hd__and2_1 c233 (.A(net157),
    .B(net197),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_1 c234 (.A(net755),
    .X(net209));
 sky130_fd_sc_hd__and2_1 c235 (.A(net18),
    .B(net171),
    .X(net210));
 sky130_fd_sc_hd__dlymetal6s2s_1 c236 (.A(net754),
    .X(net211));
 sky130_fd_sc_hd__mux4_2 c237 (.A0(net171),
    .A1(net158),
    .A2(net81),
    .A3(net210),
    .S0(net182),
    .S1(net992),
    .X(net968));
 sky130_fd_sc_hd__and2_0 c238 (.A(net210),
    .B(clknet_1_0__leaf_net855),
    .X(net212));
 sky130_fd_sc_hd__a2111o_1 c239 (.A1(net199),
    .A2(net211),
    .B1(net968),
    .C1(net992),
    .D1(net205),
    .X(net213));
 sky130_fd_sc_hd__a2111o_1 c240 (.A1(net212),
    .A2(net211),
    .B1(net210),
    .C1(net69),
    .D1(net200),
    .X(net214));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(net71),
    .A1(net206),
    .A2(net61),
    .A3(net72),
    .S0(net13),
    .S1(net837),
    .X(net215));
 sky130_fd_sc_hd__and3_4 c242 (.A(net211),
    .B(net69),
    .C(net84),
    .X(net216));
 sky130_fd_sc_hd__mux4_1 c243 (.A0(net68),
    .A1(net84),
    .A2(net99),
    .A3(net206),
    .S0(net216),
    .S1(net188),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_1 c244 (.A(net734),
    .X(net218));
 sky130_fd_sc_hd__buf_1 c245 (.A(net763),
    .X(net219));
 sky130_fd_sc_hd__or4bb_1 c246 (.A(net208),
    .B(net216),
    .C_N(net1027),
    .D_N(net68),
    .X(net220));
 sky130_fd_sc_hd__or4bb_1 c247 (.A(net188),
    .B(net1024),
    .C_N(net1007),
    .D_N(clknet_1_0__leaf_net856),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_1 c248 (.A(net943),
    .X(net222));
 sky130_fd_sc_hd__mux4_1 c249 (.A0(net87),
    .A1(net1026),
    .A2(net205),
    .A3(net35),
    .S0(net211),
    .S1(net1034),
    .X(net223));
 sky130_fd_sc_hd__and2_1 c25 (.A(net951),
    .B(net957),
    .X(net0));
 sky130_fd_sc_hd__clkbuf_1 c250 (.A(net829),
    .X(net224));
 sky130_fd_sc_hd__dlymetal6s2s_1 c251 (.A(net735),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 c252 (.A(net829),
    .X(net226));
 sky130_fd_sc_hd__sdfrtn_1 c253 (.CLK_N(clknet_4_10_0_clk),
    .D(net101),
    .RESET_B(net96),
    .SCD(net216),
    .SCE(net1007),
    .Q(net227));
 sky130_fd_sc_hd__a2111o_1 c254 (.A1(net84),
    .A2(net188),
    .B1(net114),
    .C1(net227),
    .D1(net992),
    .X(net228));
 sky130_fd_sc_hd__sdfrtp_4 c255 (.CLK(clknet_4_10_0_clk),
    .D(net228),
    .RESET_B(net227),
    .SCD(net968),
    .SCE(net1034),
    .Q(net229));
 sky130_fd_sc_hd__sdfbbp_1 c256 (.CLK(clknet_4_11_0_clk),
    .D(net158),
    .RESET_B(net104),
    .SCD(net1063),
    .SCE(net93),
    .SET_B(net96),
    .Q(net971),
    .Q_N(net230));
 sky130_fd_sc_hd__mux4_1 c257 (.A0(net226),
    .A1(net223),
    .A2(net208),
    .A3(net84),
    .S0(clknet_1_0__leaf_net221),
    .S1(net216),
    .X(net231));
 sky130_fd_sc_hd__mux4_1 c258 (.A0(net87),
    .A1(net227),
    .A2(net216),
    .A3(net99),
    .S0(net220),
    .X(net232));
 sky130_fd_sc_hd__sdfbbn_1 c259 (.CLK_N(clknet_4_11_0_clk),
    .D(net172),
    .RESET_B(net99),
    .SCD(net68),
    .SCE(net48),
    .SET_B(net96),
    .Q(net234),
    .Q_N(net233));
 sky130_fd_sc_hd__and2_4 c26 (.A(net950),
    .B(net964),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 c260 (.A(net762),
    .X(net235));
 sky130_fd_sc_hd__and3_1 c261 (.A(net235),
    .B(net227),
    .C(net234),
    .X(net236));
 sky130_fd_sc_hd__a2111o_4 c262 (.A1(net218),
    .A2(net235),
    .B1(net997),
    .C1(net813),
    .D1(net998),
    .X(net237));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net234),
    .A1(net236),
    .A2(net235),
    .A3(net68),
    .S0(net1029),
    .S1(net216),
    .X(net238));
 sky130_fd_sc_hd__and2_1 c264 (.A(net110),
    .B(net953),
    .X(net239));
 sky130_fd_sc_hd__and2_0 c265 (.A(net110),
    .B(net111),
    .X(net240));
 sky130_fd_sc_hd__and2_1 c266 (.A(net120),
    .B(net123),
    .X(net241));
 sky130_fd_sc_hd__and2_4 c267 (.A(net955),
    .B(net954),
    .X(net242));
 sky130_fd_sc_hd__and2_0 c268 (.A(net785),
    .B(net119),
    .X(net243));
 sky130_fd_sc_hd__and2_1 c269 (.A(net105),
    .B(net243),
    .X(net244));
 sky130_fd_sc_hd__and2_4 c27 (.A(net1),
    .B(net961),
    .X(net2));
 sky130_fd_sc_hd__and2_2 c270 (.A(net244),
    .B(net363),
    .X(net245));
 sky130_fd_sc_hd__and2_1 c271 (.A(net960),
    .B(net242),
    .X(net246));
 sky130_fd_sc_hd__and2_0 c272 (.A(net945),
    .B(net122),
    .X(net247));
 sky130_fd_sc_hd__and2_1 c273 (.A(net247),
    .B(net239),
    .X(net248));
 sky130_fd_sc_hd__and2_0 c274 (.A(net243),
    .B(net246),
    .X(net249));
 sky130_fd_sc_hd__and2_0 c275 (.A(net239),
    .B(net245),
    .X(net250));
 sky130_fd_sc_hd__and3_1 c276 (.A(net118),
    .B(net244),
    .C(net239),
    .X(net251));
 sky130_fd_sc_hd__and2_1 c277 (.A(net249),
    .B(net250),
    .X(net252));
 sky130_fd_sc_hd__and3_4 c278 (.A(net251),
    .B(net252),
    .C(net250),
    .X(net253));
 sky130_fd_sc_hd__and3_1 c279 (.A(net251),
    .B(net986),
    .C(net245),
    .X(net254));
 sky130_fd_sc_hd__and2_2 c28 (.A(net955),
    .B(net949),
    .X(net3));
 sky130_fd_sc_hd__and3_1 c280 (.A(net250),
    .B(net112),
    .C(net252),
    .X(net255));
 sky130_fd_sc_hd__mux4_2 c281 (.A0(net254),
    .A1(net248),
    .A2(net249),
    .A3(net241),
    .S0(net242),
    .S1(net253),
    .X(net256));
 sky130_fd_sc_hd__or4bb_2 c282 (.A(net255),
    .B(net251),
    .C_N(net954),
    .D_N(net991),
    .X(net257));
 sky130_fd_sc_hd__mux4_1 c283 (.A0(net252),
    .A1(net247),
    .A2(net257),
    .A3(net248),
    .S0(net991),
    .S1(net242),
    .X(net258));
 sky130_fd_sc_hd__and3_1 c284 (.A(net243),
    .B(net252),
    .C(net816),
    .X(net259));
 sky130_fd_sc_hd__mux4_1 c285 (.A0(net259),
    .A1(net241),
    .A2(net244),
    .A3(net255),
    .S0(net257),
    .S1(net954),
    .X(net260));
 sky130_fd_sc_hd__and2_1 c286 (.A(net146),
    .B(net3),
    .X(net261));
 sky130_fd_sc_hd__and2_2 c287 (.A(net245),
    .B(net816),
    .X(net262));
 sky130_fd_sc_hd__or4bb_2 c288 (.A(net248),
    .B(net262),
    .C_N(net5),
    .D_N(net1020),
    .X(net263));
 sky130_fd_sc_hd__and2_1 c289 (.A(net141),
    .B(net246),
    .X(net264));
 sky130_fd_sc_hd__and2_1 c29 (.A(net958),
    .B(net956),
    .X(net4));
 sky130_fd_sc_hd__and3_1 c290 (.A(net261),
    .B(net144),
    .C(net816),
    .X(net265));
 sky130_fd_sc_hd__and3_4 c291 (.A(net124),
    .B(net130),
    .C(net262),
    .X(net266));
 sky130_fd_sc_hd__buf_1 c292 (.A(net788),
    .X(net267));
 sky130_fd_sc_hd__and3_2 c293 (.A(net147),
    .B(net146),
    .C(net13),
    .X(net268));
 sky130_fd_sc_hd__and2_4 c294 (.A(net2),
    .B(net261),
    .X(net269));
 sky130_fd_sc_hd__and3_1 c295 (.A(net965),
    .B(net144),
    .C(net269),
    .X(net270));
 sky130_fd_sc_hd__or4bb_1 c296 (.A(net107),
    .B(net265),
    .C_N(net245),
    .D_N(net269),
    .X(net271));
 sky130_fd_sc_hd__or4bb_1 c297 (.A(net246),
    .B(net271),
    .C_N(net262),
    .D_N(net253),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_2 c298 (.A(net836),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_1 c299 (.A(net836),
    .X(net274));
 sky130_fd_sc_hd__and2_2 c30 (.A(net949),
    .B(net952),
    .X(net5));
 sky130_fd_sc_hd__a2111o_1 c300 (.A1(net272),
    .A2(net270),
    .B1(net800),
    .C1(net115),
    .D1(net262),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_1 c301 (.A(net788),
    .X(net276));
 sky130_fd_sc_hd__and2_1 c302 (.A(net270),
    .B(net271),
    .X(net277));
 sky130_fd_sc_hd__a2111o_1 c303 (.A1(net246),
    .A2(net267),
    .B1(net262),
    .C1(net273),
    .D1(net789),
    .X(net278));
 sky130_fd_sc_hd__sdfrtp_1 c304 (.CLK(clknet_4_0_0_clk),
    .D(net271),
    .RESET_B(net268),
    .SCD(net277),
    .SCE(net816),
    .Q(net279));
 sky130_fd_sc_hd__mux4_2 c305 (.A0(net276),
    .A1(net261),
    .A2(net279),
    .A3(net146),
    .S0(net264),
    .S1(net816),
    .X(net280));
 sky130_fd_sc_hd__or4bb_1 c306 (.A(net128),
    .B(net277),
    .C_N(net276),
    .D_N(net279),
    .X(net281));
 sky130_fd_sc_hd__mux4_1 c307 (.A0(net265),
    .A1(net263),
    .A2(net277),
    .A3(net994),
    .S0(net267),
    .S1(net245),
    .X(net282));
 sky130_fd_sc_hd__and3_2 c308 (.A(net126),
    .B(net994),
    .C(net273),
    .X(net283));
 sky130_fd_sc_hd__and3_1 c309 (.A(net136),
    .B(net279),
    .C(net1013),
    .X(net284));
 sky130_fd_sc_hd__and3_4 c31 (.A(net2),
    .B(net951),
    .C(net1),
    .X(net6));
 sky130_fd_sc_hd__and3_2 c310 (.A(net947),
    .B(net106),
    .C(net1002),
    .X(net285));
 sky130_fd_sc_hd__buf_2 c311 (.A(net1070),
    .X(net286));
 sky130_fd_sc_hd__a2111o_2 c312 (.A1(net124),
    .A2(net136),
    .B1(net165),
    .C1(net995),
    .D1(net844),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_1 c313 (.A(net924),
    .X(net288));
 sky130_fd_sc_hd__or4bb_2 c314 (.A(net108),
    .B(net1009),
    .C_N(net996),
    .D_N(net816),
    .X(net289));
 sky130_fd_sc_hd__and3_4 c315 (.A(net169),
    .B(net28),
    .C(net286),
    .X(net975));
 sky130_fd_sc_hd__and3_1 c316 (.A(net164),
    .B(net155),
    .C(net289),
    .X(net290));
 sky130_fd_sc_hd__and3_1 c317 (.A(net154),
    .B(net283),
    .C(net279),
    .X(net291));
 sky130_fd_sc_hd__buf_1 c318 (.A(clknet_1_0__leaf_net931),
    .X(net292));
 sky130_fd_sc_hd__mux4_1 c319 (.A0(net288),
    .A1(net975),
    .A2(net136),
    .A3(net1014),
    .S0(net131),
    .S1(net144),
    .X(net293));
 sky130_fd_sc_hd__and2_1 c32 (.A(net964),
    .B(net3),
    .X(net7));
 sky130_fd_sc_hd__and3_1 c320 (.A(net279),
    .B(net245),
    .C(net144),
    .X(net294));
 sky130_fd_sc_hd__and3_1 c321 (.A(net363),
    .B(net274),
    .C(net279),
    .X(net295));
 sky130_fd_sc_hd__mux4_1 c322 (.A0(net155),
    .A1(net273),
    .A2(clknet_1_0__leaf_net292),
    .A3(net294),
    .S0(net291),
    .S1(net843),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_1 c323 (.A(net939),
    .X(net297));
 sky130_fd_sc_hd__mux4_1 c324 (.A0(net277),
    .A1(net269),
    .A2(net165),
    .A3(net287),
    .S0(net844),
    .S1(net859),
    .X(net298));
 sky130_fd_sc_hd__and3_1 c325 (.A(net844),
    .B(net860),
    .C(net862),
    .X(net299));
 sky130_fd_sc_hd__mux4_1 c326 (.A0(net294),
    .A1(net295),
    .A2(net164),
    .A3(net299),
    .S0(net253),
    .S1(net287),
    .X(net300));
 sky130_fd_sc_hd__mux4_2 c327 (.A0(net295),
    .A1(net995),
    .A2(net299),
    .A3(net994),
    .S0(net245),
    .S1(net857),
    .X(net301));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(net290),
    .A1(net294),
    .A2(net283),
    .A3(net299),
    .S0(net6),
    .S1(net860),
    .X(net302));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net115),
    .A1(net299),
    .A2(net277),
    .S0(net857),
    .S1(net863),
    .X(net303));
 sky130_fd_sc_hd__and2_4 c33 (.A(net964),
    .B(net951),
    .X(net8));
 sky130_fd_sc_hd__and2_2 c330 (.A(net151),
    .B(net816),
    .X(net304));
 sky130_fd_sc_hd__a2111o_1 c331 (.A1(net269),
    .A2(net180),
    .B1(net285),
    .C1(net304),
    .D1(clknet_1_0__leaf_net854),
    .X(net305));
 sky130_fd_sc_hd__dlymetal6s2s_1 c332 (.A(net837),
    .X(net306));
 sky130_fd_sc_hd__and2_2 c333 (.A(net8),
    .B(net306),
    .X(net307));
 sky130_fd_sc_hd__and2_0 c334 (.A(net306),
    .B(net860),
    .X(net308));
 sky130_fd_sc_hd__and3_1 c335 (.A(net55),
    .B(net39),
    .C(clknet_1_0__leaf_net854),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_1 c336 (.A(net837),
    .X(net310));
 sky130_fd_sc_hd__sdfbbn_1 c337 (.CLK_N(clknet_4_9_0_clk),
    .D(net306),
    .RESET_B(net268),
    .SCD(net191),
    .SCE(net304),
    .SET_B(net1043),
    .Q(net312),
    .Q_N(net311));
 sky130_fd_sc_hd__and2_0 c338 (.A(net816),
    .B(net863),
    .X(net313));
 sky130_fd_sc_hd__and3_1 c339 (.A(net310),
    .B(net8),
    .C(net311),
    .X(net314));
 sky130_fd_sc_hd__and2_1 c34 (.A(net4),
    .B(net6),
    .X(net9));
 sky130_fd_sc_hd__and3_1 c340 (.A(net309),
    .B(net312),
    .C(net304),
    .X(net315));
 sky130_fd_sc_hd__mux4_1 c341 (.A0(net312),
    .A1(net310),
    .A2(net306),
    .A3(net994),
    .S0(net48),
    .S1(net304),
    .X(net316));
 sky130_fd_sc_hd__mux4_1 c342 (.A0(net291),
    .A1(net289),
    .A2(net312),
    .A3(clknet_1_0__leaf_net315),
    .S0(net306),
    .S1(net304),
    .X(net317));
 sky130_fd_sc_hd__and2_0 c343 (.A(net307),
    .B(net843),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_1 c344 (.A(net777),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_2 c345 (.A(net776),
    .X(net320));
 sky130_fd_sc_hd__mux4_1 c346 (.A0(net320),
    .A1(clknet_1_0__leaf_net315),
    .A2(net318),
    .A3(net807),
    .S0(net843),
    .S1(clknet_1_0__leaf_net854),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_1 c347 (.A(net932),
    .X(net322));
 sky130_fd_sc_hd__and3_2 c348 (.A(net319),
    .B(net993),
    .C(net865),
    .X(net323));
 sky130_fd_sc_hd__and2_1 c349 (.A(net322),
    .B(net323),
    .X(net324));
 sky130_fd_sc_hd__and2_2 c35 (.A(net5),
    .B(net7),
    .X(net10));
 sky130_fd_sc_hd__or4bb_1 c350 (.A(net187),
    .B(net306),
    .C_N(net323),
    .D_N(net191),
    .X(net325));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net324),
    .A1(net311),
    .A2(net320),
    .A3(net991),
    .S0(net806),
    .S1(net857),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_1 c352 (.A(net768),
    .X(net327));
 sky130_fd_sc_hd__and2_1 c353 (.A(net114),
    .B(net864),
    .X(net328));
 sky130_fd_sc_hd__buf_1 c354 (.A(clknet_1_1__leaf_net931),
    .X(net329));
 sky130_fd_sc_hd__and2_1 c355 (.A(net327),
    .B(net800),
    .X(net330));
 sky130_fd_sc_hd__and2_0 c356 (.A(net200),
    .B(net304),
    .X(net331));
 sky130_fd_sc_hd__and2_1 c357 (.A(net209),
    .B(net78),
    .X(net332));
 sky130_fd_sc_hd__and2_0 c358 (.A(net794),
    .B(clknet_1_1__leaf_net855),
    .X(net333));
 sky130_fd_sc_hd__and2_2 c359 (.A(net198),
    .B(net200),
    .X(net334));
 sky130_fd_sc_hd__and2_4 c36 (.A(net10),
    .B(net9),
    .X(net11));
 sky130_fd_sc_hd__mux4_1 c360 (.A0(net332),
    .A1(net304),
    .A2(net998),
    .A3(clknet_1_1__leaf_net315),
    .S0(net799),
    .S1(clknet_1_1__leaf_net855),
    .X(net335));
 sky130_fd_sc_hd__and3_1 c361 (.A(net297),
    .B(net327),
    .C(clknet_1_1__leaf_net854),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_1 c362 (.A(net725),
    .X(net337));
 sky130_fd_sc_hd__and2_0 c363 (.A(clknet_1_1__leaf_net329),
    .B(net866),
    .X(net338));
 sky130_fd_sc_hd__buf_1 c364 (.A(net937),
    .X(net339));
 sky130_fd_sc_hd__mux4_2 c365 (.A0(net78),
    .A1(clknet_1_0__leaf_net329),
    .A2(net997),
    .A3(net269),
    .S0(net205),
    .S1(clknet_1_0__leaf_net823),
    .X(net985));
 sky130_fd_sc_hd__clkbuf_1 c366 (.A(net725),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_2 c367 (.A(net751),
    .X(net341));
 sky130_fd_sc_hd__or4bb_1 c368 (.A(net331),
    .B(net341),
    .C_N(net992),
    .D_N(clknet_1_1__leaf_net854),
    .X(net342));
 sky130_fd_sc_hd__and2_0 c369 (.A(net340),
    .B(clknet_1_1__leaf_net854),
    .X(net969));
 sky130_fd_sc_hd__and2_1 c37 (.A(net956),
    .B(net4),
    .X(net12));
 sky130_fd_sc_hd__mux4_1 c370 (.A0(net336),
    .A1(net200),
    .A2(clknet_1_0__leaf_net969),
    .A3(net341),
    .S0(net48),
    .S1(net334),
    .X(net343));
 sky130_fd_sc_hd__sdfrtp_1 c371 (.CLK(clknet_4_9_0_clk),
    .D(net48),
    .RESET_B(clknet_1_0__leaf_net969),
    .SCD(clknet_1_1__leaf_net854),
    .SCE(net857),
    .Q(net344));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net337),
    .A1(clknet_1_0__leaf_net969),
    .A2(clknet_1_1__leaf_net315),
    .A3(net334),
    .S0(clknet_1_0__leaf_net823),
    .S1(net867),
    .X(net345));
 sky130_fd_sc_hd__or4bb_1 c373 (.A(net341),
    .B(clknet_1_1__leaf_net823),
    .C_N(net866),
    .D_N(net868),
    .X(net346));
 sky130_fd_sc_hd__mux4_1 c374 (.A0(net206),
    .A1(net227),
    .A2(net237),
    .A3(net975),
    .S0(net191),
    .S1(net847),
    .X(net347));
 sky130_fd_sc_hd__sdfsbp_1 c375 (.CLK(clknet_4_11_0_clk),
    .D(clknet_1_1__leaf_net315),
    .SCD(net992),
    .SCE(net227),
    .SET_B(clknet_1_0__leaf_net969),
    .Q(net349),
    .Q_N(net348));
 sky130_fd_sc_hd__a2111o_1 c376 (.A1(net1030),
    .A2(net222),
    .B1(net330),
    .C1(net6),
    .D1(net1007),
    .X(net350));
 sky130_fd_sc_hd__sdfsbp_1 c377 (.CLK(clknet_4_11_0_clk),
    .D(net350),
    .SCD(net93),
    .SCE(net216),
    .SET_B(net1050),
    .Q(net352),
    .Q_N(net351));
 sky130_fd_sc_hd__a2111o_1 c378 (.A1(net216),
    .A2(net229),
    .B1(net1034),
    .C1(net853),
    .D1(clknet_1_1__leaf_net856),
    .X(net353));
 sky130_fd_sc_hd__or4bb_1 c379 (.A(net333),
    .B(net99),
    .C_N(net229),
    .D_N(net869),
    .X(net974));
 sky130_fd_sc_hd__mux4_2 c38 (.A0(net2),
    .A1(net956),
    .A2(net12),
    .A3(net6),
    .S0(net957),
    .S1(net3),
    .X(net979));
 sky130_fd_sc_hd__mux4_2 c380 (.A0(net69),
    .A1(net99),
    .A2(net219),
    .A3(clknet_1_0__leaf_net974),
    .S0(net997),
    .S1(net237),
    .X(net354));
 sky130_fd_sc_hd__sdfstp_1 c381 (.CLK(clknet_4_11_0_clk),
    .D(net238),
    .SCD(net191),
    .SCE(clknet_1_0__leaf_net353),
    .SET_B(net1047),
    .Q(net355));
 sky130_fd_sc_hd__mux4_1 c382 (.A0(net48),
    .A1(net349),
    .A2(net191),
    .A3(net991),
    .S0(clknet_1_0__leaf_net354),
    .S1(net1008),
    .X(net356));
 sky130_fd_sc_hd__a2111o_1 c383 (.A1(net219),
    .A2(clknet_1_0__leaf_net353),
    .B1(net1008),
    .C1(clknet_1_1__leaf_net969),
    .D1(net93),
    .X(net357));
 sky130_fd_sc_hd__mux4_1 c384 (.A0(net352),
    .A1(net48),
    .A2(clknet_1_0__leaf_net354),
    .A3(net93),
    .S0(clknet_1_0__leaf_net856),
    .S1(net858),
    .X(net358));
 sky130_fd_sc_hd__a2111o_1 c385 (.A1(net216),
    .A2(net328),
    .B1(net93),
    .C1(net99),
    .D1(net1008),
    .X(net359));
 sky130_fd_sc_hd__sdfbbp_1 c386 (.CLK(clknet_4_14_0_clk),
    .D(net289),
    .RESET_B(net357),
    .SCD(net222),
    .SCE(clknet_1_1__leaf_net354),
    .SET_B(net1008),
    .Q(net988),
    .Q_N(net360));
 sky130_fd_sc_hd__or4bb_4 c387 (.A(net6),
    .B(clknet_1_0__leaf_net985),
    .C_N(net172),
    .D_N(net871),
    .X(net361));
 sky130_fd_sc_hd__mux4_2 c388 (.A0(net971),
    .A1(net348),
    .A2(net1008),
    .A3(net172),
    .S0(clknet_1_0__leaf_net830),
    .S1(net1007),
    .X(net362));
 sky130_fd_sc_hd__mux4_2 c389 (.A0(clknet_1_0__leaf_net361),
    .A1(net93),
    .A2(clknet_1_0__leaf_net354),
    .A3(net992),
    .S1(clknet_1_1__leaf_net856),
    .X(net830));
 sky130_fd_sc_hd__a2111o_4 c39 (.A1(net12),
    .A2(net10),
    .B1(net8),
    .C1(net11),
    .D1(net979),
    .X(net13));
 sky130_fd_sc_hd__sdfbbn_1 c390 (.CLK_N(clknet_4_11_0_clk),
    .D(net362),
    .RESET_B(net172),
    .SCD(clknet_1_1__leaf_net361),
    .SCE(net359),
    .SET_B(net1008),
    .Q(net365),
    .Q_N(net364));
 sky130_fd_sc_hd__a2111o_1 c391 (.A1(net304),
    .A2(net359),
    .B1(net360),
    .C1(net963),
    .D1(net1007),
    .X(net366));
 sky130_fd_sc_hd__sdfbbn_1 c392 (.CLK_N(clknet_4_14_0_clk),
    .D(net330),
    .RESET_B(net350),
    .SCD(clknet_1_1__leaf_net354),
    .SCE(clknet_1_0__leaf_net974),
    .SET_B(net870),
    .Q(net368),
    .Q_N(net367));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net368),
    .A1(net238),
    .A2(net269),
    .A3(net1008),
    .S0(net364),
    .S1(clknet_1_1__leaf_net830),
    .X(net369));
 sky130_fd_sc_hd__sdfbbp_1 c394 (.CLK(clknet_4_14_0_clk),
    .D(clknet_1_1__leaf_net354),
    .RESET_B(net366),
    .SCD(net1008),
    .SCE(net360),
    .SET_B(net1039),
    .Q(net371),
    .Q_N(net370));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net365),
    .A1(net366),
    .A2(net370),
    .A3(net367),
    .S0(net1062),
    .S1(net1039),
    .X(net372));
 sky130_fd_sc_hd__and2_2 c396 (.A(net986),
    .B(net991),
    .X(net373));
 sky130_fd_sc_hd__buf_1 c397 (.A(net743),
    .X(net374));
 sky130_fd_sc_hd__and2_0 c398 (.A(net948),
    .B(net125),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_1 c399 (.A(net815),
    .X(net376));
 sky130_fd_sc_hd__a2111o_2 c40 (.A1(net4),
    .A2(net12),
    .B1(net1),
    .C1(net957),
    .D1(net951),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 c400 (.A(net743),
    .X(net377));
 sky130_fd_sc_hd__and2_1 c401 (.A(net120),
    .B(net259),
    .X(net378));
 sky130_fd_sc_hd__and2_1 c402 (.A(net375),
    .B(net240),
    .X(net379));
 sky130_fd_sc_hd__and2_2 c403 (.A(net240),
    .B(net253),
    .X(net380));
 sky130_fd_sc_hd__dlymetal6s2s_1 c404 (.A(net752),
    .X(net381));
 sky130_fd_sc_hd__and2_0 c405 (.A(net377),
    .B(net375),
    .X(net382));
 sky130_fd_sc_hd__and2_1 c406 (.A(net254),
    .B(net380),
    .X(net383));
 sky130_fd_sc_hd__and2_0 c407 (.A(net382),
    .B(net253),
    .X(net384));
 sky130_fd_sc_hd__and2_1 c408 (.A(net376),
    .B(net378),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_1 c409 (.A(net759),
    .X(net386));
 sky130_fd_sc_hd__a2111o_4 c41 (.A1(net13),
    .A2(net979),
    .B1(net14),
    .C1(net0),
    .D1(net7),
    .X(net15));
 sky130_fd_sc_hd__buf_1 c410 (.A(net759),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_2 c411 (.A(net815),
    .X(net388));
 sky130_fd_sc_hd__and2_2 c412 (.A(net386),
    .B(net382),
    .X(net389));
 sky130_fd_sc_hd__buf_1 c413 (.A(net815),
    .X(net390));
 sky130_fd_sc_hd__and3_1 c414 (.A(net384),
    .B(net388),
    .C(net389),
    .X(net391));
 sky130_fd_sc_hd__buf_2 c415 (.A(net939),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_4 c416 (.A(net846),
    .X(net984));
 sky130_fd_sc_hd__mux4_1 c417 (.A0(net379),
    .A1(net254),
    .A2(net390),
    .A3(net392),
    .S0(net380),
    .S1(net118),
    .X(net393));
 sky130_fd_sc_hd__and2_1 c418 (.A(net390),
    .B(net392),
    .X(net394));
 sky130_fd_sc_hd__and2_1 c419 (.A(net244),
    .B(net266),
    .X(net395));
 sky130_fd_sc_hd__mux4_2 c42 (.A0(net9),
    .A1(net15),
    .A2(net13),
    .A3(net961),
    .S0(net8),
    .S1(net14),
    .X(net16));
 sky130_fd_sc_hd__and2_1 c420 (.A(net267),
    .B(net262),
    .X(net396));
 sky130_fd_sc_hd__and2_1 c421 (.A(net379),
    .B(net242),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_1 c422 (.A(net798),
    .X(net398));
 sky130_fd_sc_hd__and3_1 c423 (.A(net131),
    .B(net986),
    .C(net396),
    .X(net399));
 sky130_fd_sc_hd__and3_1 c424 (.A(net387),
    .B(net390),
    .C(net130),
    .X(net400));
 sky130_fd_sc_hd__and3_1 c425 (.A(net130),
    .B(net396),
    .C(net994),
    .X(net401));
 sky130_fd_sc_hd__and3_2 c426 (.A(net401),
    .B(net400),
    .C(net269),
    .X(net402));
 sky130_fd_sc_hd__and2_1 c427 (.A(net398),
    .B(net394),
    .X(net403));
 sky130_fd_sc_hd__and3_1 c428 (.A(net398),
    .B(net273),
    .C(net266),
    .X(net404));
 sky130_fd_sc_hd__and2_1 c429 (.A(net278),
    .B(net267),
    .X(net405));
 sky130_fd_sc_hd__mux4_2 c43 (.A0(net15),
    .A1(net955),
    .A2(net7),
    .A3(net14),
    .S0(net9),
    .S1(net16),
    .X(net17));
 sky130_fd_sc_hd__and3_1 c430 (.A(net397),
    .B(net396),
    .C(net399),
    .X(net406));
 sky130_fd_sc_hd__buf_1 c431 (.A(net798),
    .X(net407));
 sky130_fd_sc_hd__sdfstp_1 c432 (.CLK(clknet_4_1_0_clk),
    .D(net399),
    .SCD(net131),
    .SCE(net1019),
    .SET_B(net402),
    .Q(net408));
 sky130_fd_sc_hd__and3_1 c433 (.A(net5),
    .B(net404),
    .C(net381),
    .X(net409));
 sky130_fd_sc_hd__and3_1 c434 (.A(net396),
    .B(net388),
    .C(net405),
    .X(net410));
 sky130_fd_sc_hd__and3_1 c435 (.A(net400),
    .B(net409),
    .C(net405),
    .X(net411));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net405),
    .A1(net262),
    .A2(net402),
    .A3(net408),
    .S0(net395),
    .S1(net1021),
    .X(net412));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(net408),
    .A1(net401),
    .A2(net410),
    .A3(net407),
    .S0(net389),
    .S1(net411),
    .X(net413));
 sky130_fd_sc_hd__buf_2 c438 (.A(net797),
    .X(net414));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net404),
    .A1(net408),
    .A2(net397),
    .A3(net130),
    .S0(net392),
    .S1(net1006),
    .X(net415));
 sky130_fd_sc_hd__and2_1 c44 (.A(net16),
    .B(net6),
    .X(net18));
 sky130_fd_sc_hd__and3_1 c440 (.A(net399),
    .B(net953),
    .C(net285),
    .X(net416));
 sky130_fd_sc_hd__and3_1 c441 (.A(net263),
    .B(net407),
    .C(net283),
    .X(net417));
 sky130_fd_sc_hd__buf_1 c442 (.A(net732),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_1 c443 (.A(net731),
    .X(net419));
 sky130_fd_sc_hd__mux4_1 c444 (.A0(net418),
    .A1(net419),
    .A2(net948),
    .A3(net1002),
    .S0(net858),
    .S1(clknet_1_1__leaf_net875),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_4 c445 (.A(net941),
    .X(net421));
 sky130_fd_sc_hd__buf_1 c446 (.A(clknet_1_0__leaf_net929),
    .X(net422));
 sky130_fd_sc_hd__buf_1 c447 (.A(net933),
    .X(net423));
 sky130_fd_sc_hd__and3_1 c448 (.A(net416),
    .B(clknet_1_0__leaf_net420),
    .C(net862),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_2 c449 (.A(net944),
    .X(net425));
 sky130_fd_sc_hd__and2_1 c45 (.A(net954),
    .B(net16),
    .X(net19));
 sky130_fd_sc_hd__mux4_1 c450 (.A0(net423),
    .A1(net1002),
    .A2(net407),
    .A3(net418),
    .S0(net301),
    .S1(net421),
    .X(net426));
 sky130_fd_sc_hd__and3_1 c451 (.A(clknet_1_1__leaf_net292),
    .B(net162),
    .C(net425),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_1 c452 (.A(net941),
    .X(net428));
 sky130_fd_sc_hd__mux4_1 c453 (.A0(net395),
    .A1(net286),
    .A2(net423),
    .A3(net402),
    .S0(net421),
    .S1(clknet_1_0__leaf_net427),
    .X(net429));
 sky130_fd_sc_hd__mux4_2 c454 (.A0(net428),
    .A1(net425),
    .A2(net421),
    .A3(net423),
    .S0(net418),
    .S1(net814),
    .X(net430));
 sky130_fd_sc_hd__or4bb_1 c455 (.A(net411),
    .B(net287),
    .C_N(clknet_1_1__leaf_net424),
    .D_N(clknet_1_0__leaf_net427),
    .X(net431));
 sky130_fd_sc_hd__and3_1 c456 (.A(net299),
    .B(net421),
    .C(net814),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_1 c457 (.A(net769),
    .X(net433));
 sky130_fd_sc_hd__and3_1 c458 (.A(net433),
    .B(net430),
    .C(net425),
    .X(net434));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net430),
    .A1(clknet_1_1__leaf_net424),
    .A2(net423),
    .A3(net131),
    .S0(clknet_1_0__leaf_net427),
    .S1(clknet_1_0__leaf_net875),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_1 c46 (.A(net953),
    .X(net20));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net434),
    .A1(net283),
    .A2(net299),
    .A3(net423),
    .S0(net425),
    .S1(clknet_1_0__leaf_net876),
    .X(net436));
 sky130_fd_sc_hd__sdfbbn_2 c461 (.CLK_N(clknet_4_3_0_clk),
    .D(net422),
    .RESET_B(net287),
    .SCD(net430),
    .SCE(net857),
    .SET_B(clknet_1_1__leaf_net876),
    .Q(net438),
    .Q_N(net437));
 sky130_fd_sc_hd__or4bb_1 c462 (.A(net11),
    .B(net285),
    .C_N(net407),
    .D_N(net993),
    .X(net439));
 sky130_fd_sc_hd__or4bb_1 c463 (.A(net308),
    .B(net975),
    .C_N(net430),
    .D_N(clknet_1_1__leaf_net427),
    .X(net440));
 sky130_fd_sc_hd__and2_1 c464 (.A(net37),
    .B(net320),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_1 c465 (.A(net801),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_1 c466 (.A(net801),
    .X(net443));
 sky130_fd_sc_hd__and3_1 c467 (.A(net387),
    .B(net323),
    .C(net801),
    .X(net444));
 sky130_fd_sc_hd__and2_1 c468 (.A(net318),
    .B(net1012),
    .X(net445));
 sky130_fd_sc_hd__and3_1 c469 (.A(net961),
    .B(net242),
    .C(net984),
    .X(net446));
 sky130_fd_sc_hd__and2_1 c47 (.A(net957),
    .B(net13),
    .X(net21));
 sky130_fd_sc_hd__buf_1 c470 (.A(clknet_1_1__leaf_net929),
    .X(net447));
 sky130_fd_sc_hd__buf_1 c471 (.A(clknet_1_1__leaf_net930),
    .X(net448));
 sky130_fd_sc_hd__and2_0 c472 (.A(net443),
    .B(clknet_1_0__leaf_net448),
    .X(net449));
 sky130_fd_sc_hd__sdfstp_1 c473 (.CLK(clknet_4_9_0_clk),
    .D(net268),
    .SCD(net445),
    .SCE(net323),
    .SET_B(net191),
    .Q(net450));
 sky130_fd_sc_hd__buf_1 c474 (.A(clknet_1_0__leaf_net930),
    .X(net451));
 sky130_fd_sc_hd__and2_0 c475 (.A(clknet_1_0__leaf_net449),
    .B(net314),
    .X(net452));
 sky130_fd_sc_hd__and3_2 c476 (.A(net320),
    .B(net446),
    .C(net392),
    .X(net981));
 sky130_fd_sc_hd__mux4_2 c477 (.A0(net407),
    .A1(net392),
    .A2(net1003),
    .A3(net182),
    .S0(net960),
    .S1(net865),
    .X(net453));
 sky130_fd_sc_hd__and3_1 c478 (.A(net450),
    .B(net441),
    .C(net446),
    .X(net454));
 sky130_fd_sc_hd__or4bb_1 c479 (.A(net245),
    .B(clknet_1_0__leaf_net451),
    .C_N(clknet_1_0__leaf_net447),
    .D_N(net414),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_1 c48 (.A(net7),
    .X(net22));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net454),
    .A1(net450),
    .A2(net453),
    .A3(net1003),
    .S0(clknet_1_1__leaf_net436),
    .S1(clknet_1_0__leaf_net448),
    .X(net456));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net314),
    .A1(net994),
    .A2(net993),
    .A3(net443),
    .S0(clknet_1_1__leaf_net449),
    .S1(net323),
    .X(net457));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(net455),
    .A1(clknet_1_0__leaf_net449),
    .A2(clknet_1_0__leaf_net452),
    .A3(net1003),
    .S0(net450),
    .S1(clknet_1_0__leaf_net877),
    .X(net458));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net285),
    .A1(clknet_1_0__leaf_net458),
    .A2(net439),
    .A3(net1003),
    .S0(net848),
    .S1(clknet_1_1__leaf_net877),
    .X(net459));
 sky130_fd_sc_hd__and3_1 c484 (.A(net446),
    .B(net1001),
    .C(net203),
    .X(net460));
 sky130_fd_sc_hd__and3_1 c485 (.A(net460),
    .B(net344),
    .C(net867),
    .X(net461));
 sky130_fd_sc_hd__and3_1 c486 (.A(net963),
    .B(net341),
    .C(net421),
    .X(net462));
 sky130_fd_sc_hd__a2111o_1 c487 (.A1(net73),
    .A2(net172),
    .B1(clknet_1_0__leaf_net452),
    .C1(net51),
    .D1(net991),
    .X(net463));
 sky130_fd_sc_hd__and3_1 c488 (.A(net344),
    .B(clknet_1_0__leaf_net420),
    .C(net948),
    .X(net464));
 sky130_fd_sc_hd__a2111o_1 c489 (.A1(net203),
    .A2(net462),
    .B1(clknet_1_1__leaf_net447),
    .C1(net182),
    .D1(net334),
    .X(net465));
 sky130_fd_sc_hd__and2_1 c49 (.A(net38),
    .B(net10),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 c490 (.A(net926),
    .X(net466));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(net51),
    .A1(net460),
    .A2(net466),
    .A3(net984),
    .S0(net1002),
    .S1(net865),
    .X(net467));
 sky130_fd_sc_hd__buf_2 c492 (.A(net926),
    .X(net468));
 sky130_fd_sc_hd__and3_1 c493 (.A(net339),
    .B(net334),
    .C(net466),
    .X(net469));
 sky130_fd_sc_hd__and3_1 c494 (.A(net107),
    .B(net469),
    .C(net162),
    .X(net470));
 sky130_fd_sc_hd__or4bb_1 c495 (.A(clknet_1_0__leaf_net458),
    .B(net975),
    .C_N(net785),
    .D_N(net865),
    .X(net471));
 sky130_fd_sc_hd__clkbuf_2 c496 (.A(net750),
    .X(net472));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net462),
    .A1(clknet_1_1__leaf_net458),
    .A2(net472),
    .A3(clknet_1_0__leaf_net338),
    .S0(clknet_1_0__leaf_net463),
    .S1(net11),
    .X(net473));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(clknet_1_0__leaf_net463),
    .A1(net460),
    .A2(net472),
    .A3(net334),
    .S0(net172),
    .X(net474));
 sky130_fd_sc_hd__or4bb_1 c499 (.A(net461),
    .B(net182),
    .C_N(net472),
    .D_N(net879),
    .X(net475));
 sky130_fd_sc_hd__and2_1 c50 (.A(net22),
    .B(net21),
    .X(net24));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(net470),
    .A1(net984),
    .A2(clknet_1_0__leaf_net464),
    .A3(net1006),
    .S0(clknet_1_1__leaf_net877),
    .S1(net879),
    .X(net476));
 sky130_fd_sc_hd__and3_1 c501 (.A(clknet_1_1__leaf_net338),
    .B(net472),
    .C(net878),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(clknet_1_1__leaf_net451),
    .A1(net472),
    .A2(net469),
    .A3(clknet_1_0__leaf_net346),
    .S0(net795),
    .S1(net878),
    .X(net478));
 sky130_fd_sc_hd__sdfbbn_1 c503 (.CLK_N(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net464),
    .RESET_B(net1067),
    .SCD(net253),
    .SCE(net1006),
    .SET_B(net475),
    .Q(net480),
    .Q_N(net479));
 sky130_fd_sc_hd__or4bb_1 c504 (.A(clknet_1_1__leaf_net447),
    .B(net478),
    .C_N(net480),
    .D_N(net1003),
    .X(net481));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(clknet_1_1__leaf_net346),
    .A1(clknet_1_1__leaf_net464),
    .A2(clknet_1_0__leaf_net481),
    .A3(net479),
    .S0(clknet_1_1__leaf_net463),
    .S1(net839),
    .X(net482));
 sky130_fd_sc_hd__a2111o_1 c509 (.A1(net355),
    .A2(net269),
    .B1(clknet_1_0__leaf_net969),
    .C1(net472),
    .D1(net858),
    .X(net483));
 sky130_fd_sc_hd__and3_2 c51 (.A(net21),
    .B(net946),
    .C(net38),
    .X(net25));
 sky130_fd_sc_hd__a2111o_1 c510 (.A1(net328),
    .A2(net201),
    .B1(net370),
    .C1(net93),
    .D1(net1007),
    .X(net484));
 sky130_fd_sc_hd__a2111o_1 c511 (.A1(net1002),
    .A2(net93),
    .B1(net1008),
    .C1(net873),
    .D1(net881),
    .X(net485));
 sky130_fd_sc_hd__a2111o_1 c512 (.A1(net229),
    .A2(net485),
    .B1(net162),
    .C1(net114),
    .D1(net848),
    .X(net486));
 sky130_fd_sc_hd__mux4_1 c513 (.A0(net93),
    .A1(net224),
    .A2(net360),
    .A3(net1008),
    .S0(net225),
    .S1(net873),
    .X(net487));
 sky130_fd_sc_hd__mux4_1 c514 (.A0(clknet_1_1__leaf_net221),
    .A1(net486),
    .A2(net988),
    .A3(clknet_1_0__leaf_net974),
    .S0(net992),
    .S1(net1007),
    .X(net488));
 sky130_fd_sc_hd__sdfbbp_1 c515 (.CLK(clknet_4_14_0_clk),
    .D(net968),
    .RESET_B(net1052),
    .SCD(clknet_1_1__leaf_net974),
    .SCE(net1055),
    .SET_B(net1045),
    .Q(net977),
    .Q_N(net489));
 sky130_fd_sc_hd__mux4_1 c516 (.A0(net371),
    .A1(net487),
    .A2(net968),
    .A3(net1003),
    .S0(net162),
    .S1(net466),
    .X(net490));
 sky130_fd_sc_hd__a2111o_1 c517 (.A1(net81),
    .A2(net477),
    .B1(clknet_1_1__leaf_net353),
    .C1(clknet_1_1__leaf_net452),
    .D1(net229),
    .X(net983));
 sky130_fd_sc_hd__mux4_1 c518 (.A0(net981),
    .A1(net225),
    .A2(net485),
    .A3(net466),
    .S0(clknet_1_0__leaf_net983),
    .S1(net883),
    .X(net491));
 sky130_fd_sc_hd__a2111o_1 c519 (.A1(net483),
    .A2(clknet_1_1__leaf_net353),
    .B1(net988),
    .C1(clknet_1_1__leaf_net983),
    .D1(net191),
    .X(net492));
 sky130_fd_sc_hd__and2_0 c52 (.A(net1002),
    .B(net22),
    .X(net26));
 sky130_fd_sc_hd__a2111o_1 c520 (.A1(net225),
    .A2(net119),
    .B1(clknet_1_0__leaf_net974),
    .C1(net355),
    .D1(clknet_1_0__leaf_net983),
    .X(net493));
 sky130_fd_sc_hd__sdfbbn_1 c521 (.CLK_N(clknet_4_14_0_clk),
    .D(clknet_1_1__leaf_net452),
    .RESET_B(net998),
    .SCD(net963),
    .SCE(net988),
    .SET_B(clknet_1_1__leaf_net983),
    .Q(net494));
 sky130_fd_sc_hd__sdfbbn_1 c522 (.CLK_N(clknet_4_15_0_clk),
    .D(net466),
    .RESET_B(net489),
    .SCD(clknet_1_0__leaf_net983),
    .SCE(net810),
    .SET_B(net1048),
    .Q(net987));
 sky130_fd_sc_hd__mux4_1 c523 (.A0(net441),
    .A1(net484),
    .A2(net977),
    .A3(net229),
    .S0(clknet_1_1__leaf_net983),
    .S1(net880),
    .X(net495));
 sky130_fd_sc_hd__a2111o_1 c524 (.A1(net466),
    .A2(clknet_1_0__leaf_net983),
    .B1(net992),
    .C1(net811),
    .D1(net883),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c525 (.A0(net472),
    .A1(net494),
    .A2(net8),
    .A3(clknet_1_1__leaf_net983),
    .S0(net873),
    .S1(net882),
    .X(net497));
 sky130_fd_sc_hd__a2111o_1 c526 (.A1(net324),
    .A2(net475),
    .B1(net371),
    .C1(clknet_1_0__leaf_net983),
    .D1(net982),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c527 (.A0(net119),
    .A1(clknet_1_0__leaf_net974),
    .A2(clknet_1_0__leaf_net983),
    .A3(net841),
    .S0(net966),
    .S1(net982),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_4 c528 (.A(net796),
    .X(net500));
 sky130_fd_sc_hd__and2_2 c529 (.A(net259),
    .B(net500),
    .X(net501));
 sky130_fd_sc_hd__and2_1 c53 (.A(net24),
    .B(net23),
    .X(net27));
 sky130_fd_sc_hd__and2_0 c530 (.A(net947),
    .B(net501),
    .X(net502));
 sky130_fd_sc_hd__and2_1 c531 (.A(net111),
    .B(net500),
    .X(net503));
 sky130_fd_sc_hd__and2_1 c532 (.A(net386),
    .B(net377),
    .X(net504));
 sky130_fd_sc_hd__and3_1 c533 (.A(net117),
    .B(net392),
    .C(net963),
    .X(net505));
 sky130_fd_sc_hd__and2_0 c534 (.A(net125),
    .B(net253),
    .X(net506));
 sky130_fd_sc_hd__and2_1 c535 (.A(net505),
    .B(net984),
    .X(net507));
 sky130_fd_sc_hd__and2_2 c536 (.A(net253),
    .B(net125),
    .X(net508));
 sky130_fd_sc_hd__and2_0 c537 (.A(net505),
    .B(net508),
    .X(net509));
 sky130_fd_sc_hd__and2_0 c538 (.A(net508),
    .B(net380),
    .X(net510));
 sky130_fd_sc_hd__and2_1 c539 (.A(net501),
    .B(net506),
    .X(net511));
 sky130_fd_sc_hd__and3_2 c54 (.A(net24),
    .B(net26),
    .C(net1002),
    .X(net28));
 sky130_fd_sc_hd__and2_1 c540 (.A(net506),
    .B(net503),
    .X(net512));
 sky130_fd_sc_hd__clkbuf_1 c541 (.A(net796),
    .X(net513));
 sky130_fd_sc_hd__clkbuf_1 c542 (.A(net796),
    .X(net514));
 sky130_fd_sc_hd__clkbuf_1 c543 (.A(net796),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c544 (.A0(net514),
    .A1(net501),
    .A2(net952),
    .A3(net509),
    .S0(net504),
    .S1(net508),
    .X(net516));
 sky130_fd_sc_hd__and2_0 c545 (.A(net504),
    .B(net513),
    .X(net517));
 sky130_fd_sc_hd__and2_1 c546 (.A(net113),
    .B(net517),
    .X(net518));
 sky130_fd_sc_hd__clkbuf_2 c547 (.A(net758),
    .X(net519));
 sky130_fd_sc_hd__or4bb_1 c548 (.A(net513),
    .B(net519),
    .C_N(net505),
    .D_N(net884),
    .X(net520));
 sky130_fd_sc_hd__and2_1 c549 (.A(net520),
    .B(net515),
    .X(net521));
 sky130_fd_sc_hd__and2_0 c55 (.A(net960),
    .B(net1002),
    .X(net29));
 sky130_fd_sc_hd__and2_2 c550 (.A(net956),
    .B(net874),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 c551 (.A0(net394),
    .A1(net519),
    .A2(net415),
    .A3(net396),
    .S0(net501),
    .S1(net273),
    .X(net523));
 sky130_fd_sc_hd__and3_1 c552 (.A(net374),
    .B(net508),
    .C(net1006),
    .X(net524));
 sky130_fd_sc_hd__and3_1 c553 (.A(net409),
    .B(net994),
    .C(net396),
    .X(net525));
 sky130_fd_sc_hd__and2_0 c554 (.A(net263),
    .B(net273),
    .X(net526));
 sky130_fd_sc_hd__clkbuf_1 c555 (.A(net809),
    .X(net527));
 sky130_fd_sc_hd__and3_4 c556 (.A(net526),
    .B(net518),
    .C(net522),
    .X(net976));
 sky130_fd_sc_hd__and2_0 c557 (.A(net396),
    .B(net394),
    .X(net528));
 sky130_fd_sc_hd__buf_1 c558 (.A(net808),
    .X(net529));
 sky130_fd_sc_hd__clkbuf_1 c559 (.A(net1054),
    .X(net530));
 sky130_fd_sc_hd__and2_0 c56 (.A(net26),
    .B(net29),
    .X(net30));
 sky130_fd_sc_hd__buf_1 c560 (.A(net846),
    .X(net531));
 sky130_fd_sc_hd__clkbuf_1 c561 (.A(net846),
    .X(net532));
 sky130_fd_sc_hd__and2_1 c562 (.A(net528),
    .B(net507),
    .X(net533));
 sky130_fd_sc_hd__and3_1 c563 (.A(net527),
    .B(net530),
    .C(net531),
    .X(net534));
 sky130_fd_sc_hd__and2_0 c564 (.A(net378),
    .B(net533),
    .X(net535));
 sky130_fd_sc_hd__clkbuf_1 c565 (.A(net815),
    .X(net536));
 sky130_fd_sc_hd__and2_1 c566 (.A(net501),
    .B(net381),
    .X(net537));
 sky130_fd_sc_hd__clkbuf_4 c567 (.A(net935),
    .X(net538));
 sky130_fd_sc_hd__mux4_1 c568 (.A0(net534),
    .A1(net512),
    .A2(net537),
    .A3(net508),
    .S0(net976),
    .S1(net1056),
    .X(net539));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(net262),
    .A1(net536),
    .A2(net537),
    .A3(net538),
    .S0(net521),
    .S1(net886),
    .X(net540));
 sky130_fd_sc_hd__and2_2 c57 (.A(net20),
    .B(net0),
    .X(net31));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net415),
    .A1(net531),
    .A2(net537),
    .A3(net266),
    .S0(net538),
    .S1(net886),
    .X(net541));
 sky130_fd_sc_hd__mux4_1 c571 (.A0(net3),
    .A1(net537),
    .A2(net406),
    .A3(net885),
    .S0(net887),
    .S1(net1065),
    .X(net542));
 sky130_fd_sc_hd__and3_1 c572 (.A(net529),
    .B(net522),
    .C(net508),
    .X(net543));
 sky130_fd_sc_hd__mux4_1 c573 (.A0(net112),
    .A1(net286),
    .A2(net543),
    .A3(net421),
    .S0(clknet_1_0__leaf_net427),
    .S1(net991),
    .X(net544));
 sky130_fd_sc_hd__or4bb_1 c574 (.A(net153),
    .B(net1019),
    .C_N(clknet_1_0__leaf_net821),
    .D_N(net885),
    .X(net545));
 sky130_fd_sc_hd__and3_1 c575 (.A(net545),
    .B(net991),
    .C(net380),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_1 c576 (.A(net928),
    .X(net547));
 sky130_fd_sc_hd__sedfxbp_1 c577 (.CLK(clknet_4_6_0_clk),
    .D(net301),
    .DE(net266),
    .SCD(net512),
    .SCE(net529),
    .Q(net990),
    .Q_N(net548));
 sky130_fd_sc_hd__mux4_1 c578 (.A0(net532),
    .A1(net438),
    .A2(net119),
    .A3(net529),
    .S0(clknet_1_0__leaf_net436),
    .S1(net402),
    .X(net549));
 sky130_fd_sc_hd__clkbuf_1 c579 (.A(net928),
    .X(net550));
 sky130_fd_sc_hd__and3_4 c58 (.A(net29),
    .B(net24),
    .C(net30),
    .X(net972));
 sky130_fd_sc_hd__sedfxbp_1 c580 (.CLK(clknet_4_6_0_clk),
    .D(net381),
    .DE(net976),
    .SCD(net380),
    .SCE(clknet_1_0__leaf_net546),
    .Q(net980),
    .Q_N(net551));
 sky130_fd_sc_hd__clkbuf_1 c581 (.A(net934),
    .X(net552));
 sky130_fd_sc_hd__clkbuf_1 c582 (.A(net940),
    .X(net553));
 sky130_fd_sc_hd__clkbuf_1 c583 (.A(net940),
    .X(net554));
 sky130_fd_sc_hd__sedfxtp_1 c584 (.CLK(clknet_4_1_0_clk),
    .D(net512),
    .DE(clknet_1_0__leaf_net546),
    .SCD(net836),
    .SCE(net890),
    .Q(net555));
 sky130_fd_sc_hd__and3_1 c585 (.A(net380),
    .B(net421),
    .C(net555),
    .X(net556));
 sky130_fd_sc_hd__clkbuf_1 c586 (.A(net938),
    .X(net557));
 sky130_fd_sc_hd__and3_1 c587 (.A(net550),
    .B(net28),
    .C(net885),
    .X(net558));
 sky130_fd_sc_hd__sedfxtp_2 c588 (.CLK(clknet_4_3_0_clk),
    .D(net543),
    .DE(net999),
    .SCD(net1056),
    .SCE(net1058),
    .Q(net559));
 sky130_fd_sc_hd__sedfxtp_1 c589 (.CLK(clknet_4_6_0_clk),
    .D(net557),
    .DE(clknet_1_0__leaf_net427),
    .SCD(clknet_1_1__leaf_net420),
    .SCE(clknet_1_0__leaf_net546),
    .Q(net560));
 sky130_fd_sc_hd__and2_1 c59 (.A(net31),
    .B(net24),
    .X(net32));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(net560),
    .A1(clknet_1_0__leaf_net436),
    .A2(net11),
    .A3(net999),
    .S0(net972),
    .S1(net836),
    .X(net561));
 sky130_fd_sc_hd__or4bb_1 c591 (.A(net555),
    .B(net556),
    .C_N(net999),
    .D_N(clknet_1_0__leaf_net546),
    .X(net562));
 sky130_fd_sc_hd__or4bb_1 c592 (.A(net552),
    .B(net560),
    .C_N(net381),
    .D_N(net999),
    .X(net563));
 sky130_fd_sc_hd__sdfrbp_1 c593 (.CLK(clknet_4_6_0_clk),
    .D(net554),
    .RESET_B(net402),
    .SCD(clknet_1_1__leaf_net546),
    .SCE(net1061),
    .Q(net565),
    .Q_N(net564));
 sky130_fd_sc_hd__a2111o_1 c594 (.A1(net522),
    .A2(net508),
    .B1(net976),
    .C1(net848),
    .D1(clknet_1_0__leaf_net877),
    .X(net566));
 sky130_fd_sc_hd__a2111o_1 c595 (.A1(net430),
    .A2(net962),
    .B1(net280),
    .C1(net986),
    .D1(clknet_1_0__leaf_net877),
    .X(net567));
 sky130_fd_sc_hd__mux4_1 c596 (.A0(net442),
    .A1(net307),
    .A2(net1003),
    .A3(net999),
    .S0(net519),
    .S1(clknet_1_0__leaf_net877),
    .X(net568));
 sky130_fd_sc_hd__buf_1 c597 (.A(net927),
    .X(net569));
 sky130_fd_sc_hd__sdfbbp_1 c598 (.CLK(clknet_4_3_0_clk),
    .D(net153),
    .RESET_B(net414),
    .SCD(net1060),
    .SCE(clknet_1_0__leaf_net546),
    .SET_B(net999),
    .Q(net571),
    .Q_N(net570));
 sky130_fd_sc_hd__and3_1 c599 (.A(net519),
    .B(net389),
    .C(net307),
    .X(net572));
 sky130_fd_sc_hd__and3_1 c60 (.A(net32),
    .B(net29),
    .C(net31),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 c600 (.A(net927),
    .X(net573));
 sky130_fd_sc_hd__and3_1 c601 (.A(net507),
    .B(net538),
    .C(net573),
    .X(net574));
 sky130_fd_sc_hd__a2111o_1 c602 (.A1(net445),
    .A2(net538),
    .B1(net569),
    .C1(net573),
    .D1(net307),
    .X(net575));
 sky130_fd_sc_hd__and3_1 c603 (.A(net180),
    .B(net960),
    .C(net569),
    .X(net576));
 sky130_fd_sc_hd__or4bb_1 c604 (.A(net576),
    .B(net444),
    .C_N(net1059),
    .D_N(net570),
    .X(net577));
 sky130_fd_sc_hd__or4bb_2 c605 (.A(net575),
    .B(net307),
    .C_N(net522),
    .D_N(net892),
    .X(net578));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net547),
    .A1(net569),
    .A2(net180),
    .A3(net578),
    .S0(clknet_1_0__leaf_net436),
    .S1(net174),
    .X(net579));
 sky130_fd_sc_hd__sdfrbp_1 c607 (.CLK(clknet_4_6_0_clk),
    .D(clknet_1_1__leaf_net546),
    .RESET_B(net119),
    .SCD(net805),
    .SCE(net835),
    .Q(net581),
    .Q_N(net580));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net444),
    .A1(net576),
    .A2(net548),
    .A3(net581),
    .S0(net1018),
    .S1(net570),
    .X(net582));
 sky130_fd_sc_hd__sdfrtn_1 c609 (.CLK_N(clknet_4_6_0_clk),
    .D(net578),
    .RESET_B(net1003),
    .SCD(net538),
    .SCE(net865),
    .Q(net583));
 sky130_fd_sc_hd__and3_1 c61 (.A(net30),
    .B(net20),
    .C(net972),
    .X(net34));
 sky130_fd_sc_hd__sdfbbn_1 c610 (.CLK_N(clknet_4_6_0_clk),
    .D(net500),
    .RESET_B(net574),
    .SCD(net578),
    .SCE(net580),
    .SET_B(net573),
    .Q(net989));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net285),
    .A1(net576),
    .A2(net578),
    .A3(net994),
    .S0(net580),
    .S1(net999),
    .X(net584));
 sky130_fd_sc_hd__or4bb_1 c612 (.A(net508),
    .B(net572),
    .C_N(net576),
    .D_N(clknet_1_1__leaf_net546),
    .X(net585));
 sky130_fd_sc_hd__sdfbbn_1 c613 (.CLK_N(clknet_4_6_0_clk),
    .D(clknet_1_1__leaf_net546),
    .RESET_B(net576),
    .SCD(net538),
    .SCE(net388),
    .SET_B(net1042),
    .Q(net587),
    .Q_N(net586));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(net174),
    .A1(net421),
    .A2(net581),
    .A3(net307),
    .S0(net508),
    .S1(net809),
    .X(net588));
 sky130_fd_sc_hd__sdfbbp_1 c615 (.CLK(clknet_4_6_0_clk),
    .D(net432),
    .RESET_B(net587),
    .SCD(net578),
    .SCE(net1003),
    .SET_B(net1040),
    .Q(net590),
    .Q_N(net589));
 sky130_fd_sc_hd__sdfbbn_1 c616 (.CLK_N(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net546),
    .RESET_B(net800),
    .SCD(net968),
    .SCE(clknet_1_1__leaf_net823),
    .SET_B(net1053),
    .Q(net592),
    .Q_N(net591));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(net334),
    .A1(net467),
    .A2(net1003),
    .A3(net571),
    .S0(clknet_1_0__leaf_net481),
    .S1(net865),
    .X(net593));
 sky130_fd_sc_hd__a2111o_1 c618 (.A1(net553),
    .A2(net13),
    .B1(net591),
    .C1(net570),
    .D1(net865),
    .X(net594));
 sky130_fd_sc_hd__mux4_1 c619 (.A0(net341),
    .A1(net594),
    .A2(net571),
    .A3(net573),
    .S0(net468),
    .S1(net13),
    .X(net595));
 sky130_fd_sc_hd__or4bb_4 c62 (.A(net33),
    .B(net965),
    .C_N(net26),
    .D_N(net32),
    .X(net35));
 sky130_fd_sc_hd__sdfbbn_1 c620 (.CLK_N(clknet_4_12_0_clk),
    .D(clknet_1_0__leaf_net593),
    .RESET_B(net201),
    .SCD(net437),
    .SCE(clknet_1_1__leaf_net821),
    .SET_B(clknet_1_1__leaf_net877),
    .Q(net597),
    .Q_N(net596));
 sky130_fd_sc_hd__a2111o_1 c621 (.A1(net201),
    .A2(net1010),
    .B1(net174),
    .C1(net858),
    .D1(clknet_1_0__leaf_net877),
    .X(net598));
 sky130_fd_sc_hd__a2111o_1 c622 (.A1(net332),
    .A2(net256),
    .B1(net976),
    .C1(net580),
    .D1(net69),
    .X(net599));
 sky130_fd_sc_hd__a2111o_1 c623 (.A1(net28),
    .A2(net573),
    .B1(net468),
    .C1(net341),
    .D1(net174),
    .X(net600));
 sky130_fd_sc_hd__sdfbbp_1 c624 (.CLK(clknet_4_12_0_clk),
    .D(net182),
    .RESET_B(clknet_1_1__leaf_net593),
    .SCD(net467),
    .SCE(clknet_1_1__leaf_net877),
    .SET_B(net890),
    .Q(net602),
    .Q_N(net601));
 sky130_fd_sc_hd__a2111o_2 c625 (.A1(net592),
    .A2(net69),
    .B1(net596),
    .C1(net341),
    .D1(net847),
    .X(net603));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net388),
    .A1(clknet_1_1__leaf_net436),
    .A2(net603),
    .A3(net307),
    .S0(net792),
    .S1(clknet_1_1__leaf_net877),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(net568),
    .A1(net595),
    .A2(net182),
    .A3(net800),
    .S0(net573),
    .S1(net848),
    .X(net605));
 sky130_fd_sc_hd__a2111o_1 c628 (.A1(net597),
    .A2(clknet_1_0__leaf_net420),
    .B1(net468),
    .C1(net792),
    .D1(clknet_1_0__leaf_net894),
    .X(net606));
 sky130_fd_sc_hd__a2111o_1 c629 (.A1(net603),
    .A2(net468),
    .B1(net573),
    .C1(clknet_1_0__leaf_net605),
    .D1(clknet_1_0__leaf_net894),
    .X(net607));
 sky130_fd_sc_hd__mux4_2 c63 (.A0(net0),
    .A1(net32),
    .A2(net20),
    .A3(net22),
    .S0(net23),
    .S1(net1031),
    .X(net36));
 sky130_fd_sc_hd__a2111o_1 c630 (.A1(net13),
    .A2(net11),
    .B1(net602),
    .C1(net603),
    .D1(net865),
    .X(net608));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net307),
    .A1(net603),
    .A2(net414),
    .A3(net601),
    .S0(clknet_1_0__leaf_net567),
    .S1(net890),
    .X(net609));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net583),
    .A1(clknet_1_1__leaf_net436),
    .A2(net1002),
    .A3(net564),
    .S0(net603),
    .S1(net570),
    .X(net610));
 sky130_fd_sc_hd__a2111o_1 c633 (.A1(net182),
    .A2(net467),
    .B1(clknet_1_0__leaf_net605),
    .C1(net256),
    .X(net611));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net559),
    .A1(net602),
    .A2(net551),
    .A3(clknet_1_0__leaf_net605),
    .S0(net468),
    .S1(net890),
    .X(net612));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net608),
    .A1(clknet_1_0__leaf_net605),
    .A2(net602),
    .A3(net832),
    .S0(clknet_1_1__leaf_net877),
    .S1(net896),
    .X(net613));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net581),
    .A1(clknet_1_0__leaf_net609),
    .A2(clknet_1_1__leaf_net605),
    .A3(net826),
    .S0(clknet_1_1__leaf_net877),
    .S1(clknet_1_1__leaf_net894),
    .X(net614));
 sky130_fd_sc_hd__sdfbbn_1 c637 (.CLK_N(clknet_4_13_0_clk),
    .D(clknet_1_1__leaf_net609),
    .RESET_B(net601),
    .SCD(clknet_1_0__leaf_net481),
    .SCE(net1064),
    .SET_B(net898),
    .Q(net616),
    .Q_N(net615));
 sky130_fd_sc_hd__and3_2 c64 (.A(net35),
    .B(net32),
    .C(net34),
    .X(net37));
 sky130_fd_sc_hd__and2_1 c65 (.A(net0),
    .B(net14),
    .X(net38));
 sky130_fd_sc_hd__and2_2 c66 (.A(net34),
    .B(net19),
    .X(net39));
 sky130_fd_sc_hd__and2_1 c660 (.A(net121),
    .B(net963),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_1 c661 (.A(net831),
    .X(net618));
 sky130_fd_sc_hd__and2_2 c662 (.A(net617),
    .B(net618),
    .X(net619));
 sky130_fd_sc_hd__buf_1 c663 (.A(net831),
    .X(net620));
 sky130_fd_sc_hd__and2_1 c664 (.A(net991),
    .B(net125),
    .X(net621));
 sky130_fd_sc_hd__and2_1 c665 (.A(net515),
    .B(net617),
    .X(net622));
 sky130_fd_sc_hd__and2_1 c666 (.A(net392),
    .B(net620),
    .X(net623));
 sky130_fd_sc_hd__and2_1 c667 (.A(net517),
    .B(net623),
    .X(net624));
 sky130_fd_sc_hd__buf_1 c668 (.X(net625));
 sky130_fd_sc_hd__dlymetal6s2s_1 c669 (.A(net753),
    .X(net626));
 sky130_fd_sc_hd__and2_0 c67 (.A(net39),
    .B(net31),
    .X(net40));
 sky130_fd_sc_hd__and3_2 c670 (.A(net622),
    .B(net623),
    .C(net619),
    .X(net627));
 sky130_fd_sc_hd__and2_0 c671 (.A(net618),
    .B(net500),
    .X(net628));
 sky130_fd_sc_hd__clkbuf_1 c672 (.A(net780),
    .X(net629));
 sky130_fd_sc_hd__and2_0 c673 (.A(net629),
    .B(net1005),
    .X(net630));
 sky130_fd_sc_hd__and2_0 c674 (.A(net630),
    .B(net623),
    .X(net631));
 sky130_fd_sc_hd__buf_2 c675 (.A(net780),
    .X(net632));
 sky130_fd_sc_hd__or4bb_1 c676 (.A(net631),
    .B(net632),
    .C_N(net1005),
    .D_N(net621),
    .X(net633));
 sky130_fd_sc_hd__clkbuf_1 c677 (.A(net942),
    .X(net634));
 sky130_fd_sc_hd__and2_1 c678 (.A(net504),
    .B(net627),
    .X(net635));
 sky130_fd_sc_hd__a2111o_1 c679 (.A1(net635),
    .A2(net622),
    .B1(net627),
    .C1(net621),
    .X(net636));
 sky130_fd_sc_hd__and2_0 c68 (.A(net945),
    .B(net19),
    .X(net41));
 sky130_fd_sc_hd__and2_0 c680 (.A(net634),
    .B(net822),
    .X(net637));
 sky130_fd_sc_hd__clkbuf_1 c681 (.A(net758),
    .X(net638));
 sky130_fd_sc_hd__and2_1 c682 (.A(net533),
    .B(net994),
    .X(net639));
 sky130_fd_sc_hd__and2_0 c683 (.A(net1005),
    .B(net822),
    .X(net640));
 sky130_fd_sc_hd__and2_1 c684 (.A(net628),
    .B(net640),
    .X(net641));
 sky130_fd_sc_hd__and2_1 c685 (.A(net376),
    .B(net500),
    .X(net642));
 sky130_fd_sc_hd__and2_0 c686 (.A(net518),
    .B(net641),
    .X(net643));
 sky130_fd_sc_hd__sdfbbn_1 c687 (.CLK_N(clknet_4_5_0_clk),
    .D(net641),
    .RESET_B(net511),
    .SCD(net1004),
    .SCE(net619),
    .SET_B(net874),
    .Q(net645),
    .Q_N(net644));
 sky130_fd_sc_hd__mux4_1 c688 (.A0(net622),
    .A1(net538),
    .A2(net640),
    .A3(net632),
    .S0(net1006),
    .S1(net253),
    .X(net646));
 sky130_fd_sc_hd__buf_1 c689 (.A(net749),
    .X(net647));
 sky130_fd_sc_hd__and2_1 c69 (.A(net14),
    .B(net947),
    .X(net42));
 sky130_fd_sc_hd__and2_1 c690 (.A(net637),
    .B(net641),
    .X(net648));
 sky130_fd_sc_hd__and3_1 c691 (.A(net503),
    .B(net638),
    .C(net627),
    .X(net649));
 sky130_fd_sc_hd__sdfbbp_1 c692 (.CLK(clknet_4_5_0_clk),
    .D(net640),
    .RESET_B(net147),
    .SCD(net1005),
    .SCE(net638),
    .SET_B(net639),
    .Q(net651),
    .Q_N(net650));
 sky130_fd_sc_hd__mux4_2 c693 (.A0(net994),
    .A1(net645),
    .A2(net647),
    .A3(net533),
    .S0(net1006),
    .S1(net643),
    .X(net652));
 sky130_fd_sc_hd__a2111o_1 c694 (.A1(net645),
    .A2(net648),
    .B1(net652),
    .C1(net1004),
    .D1(net874),
    .X(net653));
 sky130_fd_sc_hd__a2111o_1 c695 (.A1(net991),
    .A2(net643),
    .B1(net644),
    .C1(net652),
    .D1(net641),
    .X(net654));
 sky130_fd_sc_hd__and2_0 c696 (.A(net147),
    .B(net651),
    .X(net655));
 sky130_fd_sc_hd__and2_2 c697 (.A(net655),
    .B(net651),
    .X(net656));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(net648),
    .A1(net650),
    .A2(net656),
    .A3(net500),
    .S0(net652),
    .S1(net812),
    .X(net657));
 sky130_fd_sc_hd__sdfbbn_1 c699 (.CLK_N(clknet_4_5_0_clk),
    .D(net115),
    .RESET_B(net656),
    .SCD(net652),
    .SCE(net619),
    .SET_B(net632),
    .Q(net659),
    .Q_N(net658));
 sky130_fd_sc_hd__and2_1 c70 (.A(net1031),
    .B(net39),
    .X(net43));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net641),
    .A1(net652),
    .A2(net1004),
    .A3(net656),
    .S0(net822),
    .S1(net899),
    .X(net660));
 sky130_fd_sc_hd__a2111o_1 c701 (.A1(net623),
    .A2(net627),
    .B1(net656),
    .C1(net652),
    .D1(net900),
    .X(net661));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net658),
    .A1(net656),
    .A2(net652),
    .A3(net1004),
    .S0(net899),
    .S1(net900),
    .X(net662));
 sky130_fd_sc_hd__mux4_2 c703 (.A0(net635),
    .A1(net812),
    .A2(net831),
    .A3(net899),
    .S0(net900),
    .S1(net901),
    .X(net663));
 sky130_fd_sc_hd__a2111o_1 c704 (.A1(net646),
    .A2(net663),
    .B1(net1005),
    .C1(net1004),
    .D1(net656),
    .X(net664));
 sky130_fd_sc_hd__and3_1 c705 (.A(net118),
    .B(net619),
    .C(net901),
    .X(net665));
 sky130_fd_sc_hd__a2111o_1 c706 (.A1(net648),
    .A2(net665),
    .B1(net1004),
    .C1(net627),
    .D1(net1066),
    .X(net666));
 sky130_fd_sc_hd__a2111o_1 c707 (.A1(net627),
    .A2(net430),
    .B1(net115),
    .C1(net999),
    .D1(net861),
    .X(net667));
 sky130_fd_sc_hd__and3_1 c708 (.A(net619),
    .B(net1001),
    .C(net1004),
    .X(net668));
 sky130_fd_sc_hd__a2111o_1 c709 (.A1(net543),
    .A2(net624),
    .B1(net266),
    .C1(net437),
    .D1(net647),
    .X(net669));
 sky130_fd_sc_hd__and2_1 c71 (.A(net19),
    .B(net36),
    .X(net44));
 sky130_fd_sc_hd__and3_1 c710 (.A(net656),
    .B(net1009),
    .C(net825),
    .X(net670));
 sky130_fd_sc_hd__buf_1 c711 (.A(net1041),
    .X(net671));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net659),
    .A1(net984),
    .A2(net1005),
    .A3(net670),
    .S0(net627),
    .S1(clknet_1_0__leaf_net821),
    .X(net672));
 sky130_fd_sc_hd__or4bb_1 c713 (.A(net511),
    .B(net162),
    .C_N(net1004),
    .D_N(net1006),
    .X(net673));
 sky130_fd_sc_hd__a2111o_1 c714 (.A1(net670),
    .A2(net627),
    .B1(net8),
    .C1(net115),
    .D1(net828),
    .X(net674));
 sky130_fd_sc_hd__sdfbbn_2 c715 (.CLK_N(clknet_4_5_0_clk),
    .D(net671),
    .RESET_B(net500),
    .SCD(net670),
    .SCE(net649),
    .SET_B(net824),
    .Q(net676),
    .Q_N(net675));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net666),
    .A1(net668),
    .A2(net543),
    .A3(net25),
    .S0(net675),
    .S1(net656),
    .X(net677));
 sky130_fd_sc_hd__and3_1 c717 (.A(net121),
    .B(net676),
    .C(net887),
    .X(net678));
 sky130_fd_sc_hd__or4bb_1 c718 (.A(net635),
    .B(net999),
    .C_N(net858),
    .D_N(net862),
    .X(net679));
 sky130_fd_sc_hd__and3_1 c719 (.A(net656),
    .B(net678),
    .C(net620),
    .X(net680));
 sky130_fd_sc_hd__and2_1 c72 (.A(net42),
    .B(net36),
    .X(net45));
 sky130_fd_sc_hd__a2111o_1 c720 (.A1(net649),
    .A2(net620),
    .B1(net675),
    .C1(net1004),
    .D1(net861),
    .X(net681));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net642),
    .A1(net670),
    .A2(net1069),
    .A3(net681),
    .S0(net671),
    .S1(net838),
    .X(net682));
 sky130_fd_sc_hd__a2111o_4 c722 (.A1(net620),
    .A2(net681),
    .B1(net675),
    .C1(net1000),
    .D1(net838),
    .X(net683));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net681),
    .A1(net679),
    .A2(net972),
    .A3(net683),
    .S0(net670),
    .S1(net658),
    .X(net684));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net680),
    .A1(net500),
    .A2(net242),
    .A3(net647),
    .S0(net683),
    .S1(net889),
    .X(net685));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net664),
    .A1(net632),
    .A2(net683),
    .A3(net828),
    .S0(net902),
    .S1(net903),
    .X(net686));
 sky130_fd_sc_hd__a2111o_1 c726 (.A1(net619),
    .A2(net590),
    .B1(net1001),
    .C1(net858),
    .D1(net904),
    .X(net687));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net1006),
    .A1(net39),
    .A2(net162),
    .A3(net619),
    .S0(net683),
    .S1(net632),
    .X(net688));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net962),
    .A1(net162),
    .A2(net114),
    .A3(net999),
    .S0(net652),
    .S1(net903),
    .X(net689));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(net266),
    .A1(net683),
    .A2(net500),
    .A3(net619),
    .S0(net652),
    .S1(net907),
    .X(net690));
 sky130_fd_sc_hd__and2_1 c73 (.A(net40),
    .B(net44),
    .X(net46));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net632),
    .A1(net647),
    .A2(net639),
    .A3(net663),
    .S0(net903),
    .S1(net906),
    .X(net691));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net652),
    .A1(net106),
    .A2(net1000),
    .A3(net683),
    .S0(net1005),
    .S1(clknet_1_0__leaf_net893),
    .X(net692));
 sky130_fd_sc_hd__a2111o_2 c732 (.A1(net1005),
    .A2(net538),
    .B1(net571),
    .C1(net903),
    .D1(net907),
    .X(net693));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net453),
    .A1(net563),
    .A2(net632),
    .A3(net1000),
    .S0(net676),
    .S1(net693),
    .X(net694));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(clknet_1_1__leaf_net457),
    .A1(net1000),
    .A2(net693),
    .A3(net619),
    .S0(net675),
    .S1(net907),
    .X(net695));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net1005),
    .A1(net820),
    .A2(net831),
    .A3(net908),
    .S0(net909),
    .S1(clknet_1_0__leaf_net911),
    .X(net696));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(net687),
    .A1(net663),
    .A2(net683),
    .A3(net908),
    .S0(net909),
    .S1(clknet_1_1__leaf_net911),
    .X(net697));
 sky130_fd_sc_hd__sdfbbp_1 c737 (.CLK(clknet_4_7_0_clk),
    .D(net587),
    .RESET_B(net665),
    .SCD(net688),
    .SCE(net453),
    .SET_B(net1046),
    .Q(net699),
    .Q_N(net698));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net639),
    .A1(net162),
    .A2(clknet_1_1__leaf_net420),
    .A3(net1005),
    .S0(net266),
    .S1(net908),
    .X(net700));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(net590),
    .A1(net687),
    .A2(net845),
    .A3(net857),
    .S0(net903),
    .S1(net909),
    .X(net701));
 sky130_fd_sc_hd__and3_1 c74 (.A(net41),
    .B(net10),
    .C(net39),
    .X(net47));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(net286),
    .A1(net639),
    .A2(net570),
    .A3(net693),
    .S0(net858),
    .S1(clknet_1_0__leaf_net912),
    .X(net702));
 sky130_fd_sc_hd__a2111o_1 c741 (.A1(clknet_1_1__leaf_net448),
    .A2(net701),
    .B1(net437),
    .C1(net906),
    .D1(clknet_1_0__leaf_net913),
    .X(net703));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(net688),
    .A1(net696),
    .A2(net984),
    .A3(net906),
    .S0(net910),
    .S1(clknet_1_0__leaf_net912),
    .X(net704));
 sky130_fd_sc_hd__a2111o_1 c743 (.A1(net106),
    .A2(net693),
    .B1(net589),
    .C1(net663),
    .D1(net901),
    .X(net705));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(net659),
    .A1(net563),
    .A2(net705),
    .A3(net1000),
    .S0(net626),
    .S1(net538),
    .X(net706));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(net697),
    .A1(net586),
    .A2(net909),
    .A3(clknet_1_1__leaf_net912),
    .S0(clknet_1_1__leaf_net913),
    .S1(net914),
    .X(net707));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net706),
    .A1(clknet_1_0__leaf_net707),
    .A2(net1000),
    .A3(net705),
    .S0(net907),
    .S1(clknet_1_0__leaf_net911),
    .X(net708));
 sky130_fd_sc_hd__a2111o_1 c747 (.A1(net705),
    .A2(net706),
    .B1(net909),
    .C1(clknet_1_0__leaf_net913),
    .D1(net915),
    .X(net709));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(clknet_1_1__leaf_net707),
    .A1(net571),
    .A2(net119),
    .A3(net615),
    .S0(net865),
    .S1(net890),
    .X(net710));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net253),
    .A1(net565),
    .A2(net616),
    .A3(net663),
    .S0(clknet_1_1__leaf_net605),
    .S1(net1002),
    .X(net711));
 sky130_fd_sc_hd__and2_4 c75 (.A(net34),
    .B(net47),
    .X(net48));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(net699),
    .A1(net624),
    .A2(net571),
    .A3(net890),
    .S0(net903),
    .S1(net909),
    .X(net712));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net693),
    .A1(net11),
    .A2(net676),
    .A3(clknet_1_0__leaf_net707),
    .S0(clknet_1_0__leaf_net895),
    .S1(net910),
    .X(net713));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net606),
    .A1(clknet_1_1__leaf_net463),
    .A2(net712),
    .A3(net663),
    .S0(net693),
    .S1(net858),
    .X(net714));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net676),
    .A1(clknet_1_1__leaf_net481),
    .A2(clknet_1_1__leaf_net707),
    .A3(net468),
    .S0(net905),
    .S1(net916),
    .X(net715));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net683),
    .A1(net571),
    .A2(clknet_1_1__leaf_net709),
    .A3(net960),
    .S0(clknet_1_1__leaf_net481),
    .S1(net663),
    .X(net716));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net624),
    .A1(net468),
    .A2(net698),
    .A3(clknet_1_1__leaf_net893),
    .S0(clknet_1_1__leaf_net895),
    .S1(net919),
    .X(net717));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(clknet_1_1__leaf_net567),
    .A1(clknet_1_1__leaf_net420),
    .A2(net616),
    .A3(clknet_1_1__leaf_net463),
    .S0(net414),
    .S1(net919),
    .X(net718));
 sky130_fd_sc_hd__mux4_2 c757 (.A0(net663),
    .A1(net703),
    .A2(clknet_1_1__leaf_net481),
    .A3(net468),
    .S0(net902),
    .S1(net919),
    .X(net719));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net1017),
    .A1(clknet_1_0__leaf_net719),
    .A2(clknet_1_1__leaf_net481),
    .A3(net865),
    .S0(net903),
    .S1(net917),
    .X(net720));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net438),
    .A1(clknet_1_1__leaf_net719),
    .A2(clknet_1_1__leaf_net605),
    .A3(net817),
    .S0(net890),
    .S1(net919),
    .X(net721));
 sky130_fd_sc_hd__and2_0 c76 (.A(net965),
    .B(net19),
    .X(net49));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net717),
    .A1(clknet_1_0__leaf_net709),
    .A2(clknet_1_0__leaf_net719),
    .A3(net840),
    .S0(net905),
    .S1(net920),
    .X(net722));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net676),
    .A1(net820),
    .A2(net848),
    .A3(net918),
    .S0(net921),
    .S1(net922),
    .X(net723));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(clknet_1_1__leaf_net605),
    .A1(net421),
    .A2(net723),
    .A3(clknet_1_1__leaf_net719),
    .S0(net909),
    .S1(net923),
    .X(net724));
 sky130_fd_sc_hd__and2_1 c77 (.A(net49),
    .B(net45),
    .X(net50));
 sky130_fd_sc_hd__and2_2 c78 (.A(net19),
    .B(net34),
    .X(net51));
 sky130_fd_sc_hd__or4bb_1 c79 (.A(net36),
    .B(net39),
    .C_N(net40),
    .D_N(net41),
    .X(net52));
 sky130_fd_sc_hd__and2_1 c80 (.A(net44),
    .B(net35),
    .X(net53));
 sky130_fd_sc_hd__buf_1 c81 (.A(net756),
    .X(net54));
 sky130_fd_sc_hd__and2_1 c82 (.A(net18),
    .B(net49),
    .X(net55));
 sky130_fd_sc_hd__mux4_2 c83 (.A0(net40),
    .A1(net957),
    .A2(net993),
    .A3(net1033),
    .S0(net961),
    .S1(net55),
    .X(net56));
 sky130_fd_sc_hd__mux4_1 c84 (.A0(net36),
    .A1(net993),
    .A2(net54),
    .A3(net49),
    .S0(net47),
    .S1(net56),
    .X(net57));
 sky130_fd_sc_hd__mux4_1 c85 (.A0(net54),
    .A1(net56),
    .A2(net961),
    .A3(net53),
    .S0(net34),
    .S1(net847),
    .X(net58));
 sky130_fd_sc_hd__a2111o_1 c86 (.A1(net56),
    .A2(net55),
    .B1(net54),
    .C1(net36),
    .D1(net847),
    .X(net59));
 sky130_fd_sc_hd__mux4_1 c87 (.A0(net56),
    .A1(net965),
    .A2(net43),
    .A3(net50),
    .S1(net850),
    .X(net60));
 sky130_fd_sc_hd__buf_1 c88 (.A(net730),
    .X(net61));
 sky130_fd_sc_hd__and2_1 c89 (.A(net43),
    .B(net28),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 c90 (.A(net730),
    .X(net63));
 sky130_fd_sc_hd__and2_0 c91 (.A(net63),
    .B(net993),
    .X(net64));
 sky130_fd_sc_hd__and2_0 c92 (.A(net963),
    .B(net847),
    .X(net65));
 sky130_fd_sc_hd__or4bb_1 c93 (.A(net65),
    .B(net61),
    .C_N(net50),
    .D_N(net43),
    .X(net66));
 sky130_fd_sc_hd__and2_0 c94 (.A(net972),
    .B(net993),
    .X(net67));
 sky130_fd_sc_hd__and2_2 c95 (.A(net23),
    .B(net993),
    .X(net68));
 sky130_fd_sc_hd__and2_4 c96 (.A(net10),
    .B(net63),
    .X(net69));
 sky130_fd_sc_hd__mux4_1 c97 (.A0(net65),
    .A1(net61),
    .A2(net48),
    .A3(net66),
    .S0(net31),
    .S1(net993),
    .X(net70));
 sky130_fd_sc_hd__and2_1 c98 (.A(net42),
    .B(net64),
    .X(net71));
 sky130_fd_sc_hd__sdfrbp_1 c99 (.CLK(clknet_4_8_0_clk),
    .D(net64),
    .RESET_B(net15),
    .SCD(net71),
    .SCE(net68),
    .Q(net73),
    .Q_N(net72));
 sky130_fd_sc_hd__sdfrtp_1 merge763 (.CLK(clknet_4_9_0_clk),
    .D(net191),
    .RESET_B(net74),
    .SCD(net789),
    .SCE(clknet_1_1__leaf_net855),
    .Q(net725));
 sky130_fd_sc_hd__sdfrtp_1 merge764 (.CLK(clknet_4_8_0_clk),
    .D(net66),
    .RESET_B(net157),
    .SCD(net174),
    .SCE(net992),
    .Q(net726));
 sky130_fd_sc_hd__or4bb_1 merge765 (.A(net75),
    .B(net79),
    .C_N(net15),
    .D_N(net48),
    .X(net727));
 sky130_fd_sc_hd__mux4_1 merge766 (.A0(net144),
    .A1(net277),
    .A2(net995),
    .A3(net284),
    .S0(net286),
    .S1(net166),
    .X(net728));
 sky130_fd_sc_hd__and3_1 merge767 (.A(net393),
    .B(net242),
    .C(net511),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_1 merge768 (.A(net936),
    .X(net730));
 sky130_fd_sc_hd__sdfbbn_1 merge769 (.CLK_N(clknet_4_1_0_clk),
    .D(net397),
    .RESET_B(net11),
    .SCD(net417),
    .SCE(net283),
    .SET_B(net266),
    .Q(net732),
    .Q_N(net731));
 sky130_fd_sc_hd__mux4_1 merge770 (.A0(clknet_1_1__leaf_net427),
    .A1(net1006),
    .A2(clknet_1_1__leaf_net458),
    .A3(net459),
    .S0(net465),
    .S1(net462),
    .X(net733));
 sky130_fd_sc_hd__sdfbbn_1 merge771 (.CLK_N(clknet_4_10_0_clk),
    .D(net91),
    .RESET_B(net973),
    .SCD(net217),
    .SCE(net208),
    .SET_B(net68),
    .Q(net735),
    .Q_N(net734));
 sky130_fd_sc_hd__mux4_1 merge772 (.A0(net538),
    .A1(clknet_1_0__leaf_net457),
    .A2(clknet_1_1__leaf_net448),
    .A3(net1015),
    .S0(net453),
    .S1(net522),
    .X(net736));
 sky130_fd_sc_hd__mux4_1 merge773 (.A0(net134),
    .A1(net374),
    .A2(net385),
    .A3(net402),
    .S0(net266),
    .S1(net405),
    .X(net737));
 sky130_fd_sc_hd__a2111o_1 merge774 (.A1(net287),
    .A2(net1023),
    .B1(net439),
    .C1(net320),
    .D1(clknet_1_1__leaf_net427),
    .X(net738));
 sky130_fd_sc_hd__or4bb_1 merge775 (.A(net525),
    .B(net518),
    .C_N(net273),
    .D_N(net976),
    .X(net739));
 sky130_fd_sc_hd__mux4_1 merge776 (.A0(net800),
    .A1(clknet_1_0__leaf_net427),
    .A2(clknet_1_0__leaf_net546),
    .A3(net389),
    .S0(net1022),
    .S1(net543),
    .X(net740));
 sky130_fd_sc_hd__or4bb_1 merge777 (.A(net377),
    .B(net383),
    .C_N(net952),
    .D_N(net512),
    .X(net741));
 sky130_fd_sc_hd__or4bb_1 merge778 (.A(net173),
    .B(net114),
    .C_N(net167),
    .D_N(net186),
    .X(net742));
 sky130_fd_sc_hd__buf_1 merge779 (.A(net942),
    .X(net743));
 sky130_fd_sc_hd__or4bb_1 merge780 (.A(net257),
    .B(net147),
    .C_N(net962),
    .D_N(net1057),
    .X(net744));
 sky130_fd_sc_hd__a2111o_1 merge781 (.A1(net152),
    .A2(net174),
    .B1(net286),
    .C1(net48),
    .D1(net1044),
    .X(net745));
 sky130_fd_sc_hd__mux4_1 merge782 (.A0(net323),
    .A1(clknet_1_1__leaf_net427),
    .A2(net445),
    .A3(net403),
    .S0(net975),
    .S1(net256),
    .X(net746));
 sky130_fd_sc_hd__mux4_1 merge783 (.A0(net426),
    .A1(net182),
    .A2(clknet_1_0__leaf_net447),
    .A3(net191),
    .S0(net37),
    .S1(net439),
    .X(net747));
 sky130_fd_sc_hd__or4bb_1 merge784 (.A(net509),
    .B(net389),
    .C_N(net510),
    .D_N(net112),
    .X(net748));
 sky130_fd_sc_hd__sdfrtp_1 merge785 (.CLK(clknet_4_4_0_clk),
    .D(net406),
    .RESET_B(net1068),
    .SCD(net521),
    .SCE(net525),
    .Q(net749));
 sky130_fd_sc_hd__sdfbbp_1 merge786 (.CLK(clknet_4_9_0_clk),
    .D(net207),
    .RESET_B(net28),
    .SCD(net242),
    .SCE(clknet_1_0__leaf_net464),
    .SET_B(clknet_1_0__leaf_net463),
    .Q(net751),
    .Q_N(net750));
 sky130_fd_sc_hd__sdfsbp_1 merge787 (.CLK(clknet_4_4_0_clk),
    .D(net621),
    .SCD(net619),
    .SCE(net380),
    .SET_B(net373),
    .Q(net753),
    .Q_N(net752));
 sky130_fd_sc_hd__sdfsbp_1 merge788 (.CLK(clknet_4_9_0_clk),
    .D(net61),
    .SCD(net71),
    .SCE(net207),
    .SET_B(net1038),
    .Q(net755),
    .Q_N(net754));
 sky130_fd_sc_hd__sdfstp_1 merge789 (.CLK(clknet_4_8_0_clk),
    .D(net46),
    .SCD(net993),
    .SCE(net88),
    .SET_B(net79),
    .Q(net756));
 sky130_fd_sc_hd__or4bb_1 merge790 (.A(net76),
    .B(net42),
    .C_N(net89),
    .D_N(net96),
    .X(net757));
 sky130_fd_sc_hd__sdfstp_1 merge791 (.CLK(clknet_4_5_0_clk),
    .D(net637),
    .SCD(net621),
    .SCE(net502),
    .SET_B(net503),
    .Q(net758));
 sky130_fd_sc_hd__buf_1 merge792 (.A(net846),
    .X(net759));
 sky130_fd_sc_hd__or4bb_1 merge793 (.A(net373),
    .B(net384),
    .C_N(net535),
    .D_N(net531),
    .X(net760));
 sky130_fd_sc_hd__mux4_1 merge794 (.A0(net78),
    .A1(clknet_1_0__leaf_net315),
    .A2(net165),
    .A3(net290),
    .S0(net287),
    .S1(net837),
    .X(net761));
 sky130_fd_sc_hd__sdfbbn_1 merge795 (.CLK_N(clknet_4_11_0_clk),
    .D(net1034),
    .RESET_B(net96),
    .SCD(net191),
    .SCE(net233),
    .SET_B(net813),
    .Q(net763),
    .Q_N(net762));
 sky130_fd_sc_hd__a2111o_1 merge796 (.A1(net264),
    .A2(net257),
    .B1(net141),
    .C1(net132),
    .D1(net271),
    .X(net764));
 sky130_fd_sc_hd__or4bb_1 merge797 (.A(net530),
    .B(net976),
    .C_N(net524),
    .D_N(net531),
    .X(net765));
 sky130_fd_sc_hd__sdfstp_1 merge798 (.CLK(clknet_4_10_0_clk),
    .D(net79),
    .SCD(net97),
    .SCE(net62),
    .SET_B(net31),
    .Q(net766));
 sky130_fd_sc_hd__mux4_1 merge799 (.A0(net417),
    .A1(net245),
    .A2(net283),
    .A3(net305),
    .S0(net154),
    .S1(net320),
    .X(net767));
 sky130_fd_sc_hd__sdfbbn_1 merge800 (.CLK_N(clknet_4_9_0_clk),
    .D(net417),
    .RESET_B(net74),
    .SCD(net172),
    .SCE(net81),
    .SET_B(net1049),
    .Q(net769),
    .Q_N(net768));
 sky130_fd_sc_hd__mux4_1 merge801 (.A0(net537),
    .A1(net531),
    .A2(clknet_1_0__leaf_net427),
    .A3(net500),
    .S0(net861),
    .S1(net885),
    .X(net770));
 sky130_fd_sc_hd__mux4_1 merge802 (.A0(net50),
    .A1(net77),
    .A2(net74),
    .A3(net44),
    .S0(net79),
    .S1(net69),
    .X(net771));
 sky130_fd_sc_hd__mux4_1 merge803 (.A0(net162),
    .A1(net74),
    .A2(net996),
    .A3(net52),
    .S0(net62),
    .S1(net849),
    .X(net772));
 sky130_fd_sc_hd__a2111o_1 merge804 (.A1(net374),
    .A2(net118),
    .B1(net373),
    .C1(net241),
    .D1(net379),
    .X(net773));
 sky130_fd_sc_hd__mux4_1 merge805 (.A0(net667),
    .A1(net1006),
    .A2(net670),
    .A3(net402),
    .S0(net389),
    .S1(net430),
    .X(net774));
 sky130_fd_sc_hd__mux4_1 merge806 (.A0(net166),
    .A1(net972),
    .A2(net295),
    .A3(net391),
    .S0(net373),
    .S1(net389),
    .X(net775));
 sky130_fd_sc_hd__sdfbbp_1 merge807 (.CLK(clknet_4_9_0_clk),
    .D(net313),
    .RESET_B(net311),
    .SCD(clknet_1_0__leaf_net315),
    .SCE(net863),
    .SET_B(net864),
    .Q(net777),
    .Q_N(net776));
 sky130_fd_sc_hd__mux4_1 merge808 (.A0(net552),
    .A1(clknet_1_0__leaf_net546),
    .A2(net385),
    .A3(net402),
    .S0(net511),
    .S1(net891),
    .X(net778));
 sky130_fd_sc_hd__mux4_1 merge809 (.A0(net953),
    .A1(net411),
    .A2(net399),
    .A3(net274),
    .S0(net425),
    .S1(clknet_1_0__leaf_net424),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_1 merge810 (.A(net784),
    .X(net780));
 sky130_fd_sc_hd__mux4_1 merge811 (.A0(net383),
    .A1(net632),
    .A2(net627),
    .A3(net241),
    .S0(net373),
    .S1(net113),
    .X(net781));
 sky130_fd_sc_hd__mux4_1 merge812 (.A0(clknet_1_0__leaf_net424),
    .A1(net417),
    .A2(net283),
    .A3(net95),
    .S0(net996),
    .S1(net963),
    .X(net782));
 sky130_fd_sc_hd__mux4_1 merge813 (.A0(net410),
    .A1(net411),
    .A2(net183),
    .A3(net171),
    .S0(net184),
    .S1(clknet_1_0__leaf_net875),
    .X(net783));
 sky130_fd_sc_hd__sdfbbn_1 merge814 (.CLK_N(clknet_4_4_0_clk),
    .D(net114),
    .RESET_B(net621),
    .SCD(net947),
    .SCE(net125),
    .Q(net625),
    .Q_N(net784));
 sky130_fd_sc_hd__mux4_1 merge815 (.A0(net122),
    .A1(net391),
    .A2(net390),
    .A3(net383),
    .S0(net378),
    .S1(net954),
    .X(net786));
 sky130_fd_sc_hd__mux4_1 merge816 (.A0(net220),
    .A1(net96),
    .A2(clknet_1_0__leaf_net221),
    .A3(net84),
    .S0(net819),
    .S1(net1050),
    .X(net787));
 sky130_fd_sc_hd__dfrbp_1 merge817 (.CLK(clknet_4_0_0_clk),
    .D(net275),
    .RESET_B(net744),
    .Q(net789),
    .Q_N(net788));
 sky130_fd_sc_hd__dfrbp_1 merge818 (.CLK(clknet_4_2_0_clk),
    .D(net185),
    .RESET_B(net742),
    .Q(net791),
    .Q_N(net790));
 sky130_fd_sc_hd__dfrtn_1 merge819 (.CLK_N(clknet_4_6_0_clk),
    .D(net598),
    .RESET_B(net599),
    .Q(net792));
 sky130_fd_sc_hd__and2_0 merge820 (.A(net347),
    .B(net356),
    .X(net793));
 sky130_fd_sc_hd__dfrtp_1 merge821 (.CLK(clknet_4_9_0_clk),
    .D(net204),
    .RESET_B(net214),
    .Q(net794));
 sky130_fd_sc_hd__dfrtp_1 merge822 (.CLK(clknet_4_14_0_clk),
    .D(net471),
    .Q(net474));
 sky130_fd_sc_hd__dfrtp_1 merge823 (.CLK(clknet_4_4_0_clk),
    .D(net741),
    .RESET_B(net748),
    .Q(net796));
 sky130_fd_sc_hd__dfsbp_1 merge824 (.CLK(clknet_4_0_0_clk),
    .D(net737),
    .SET_B(net783),
    .Q(net798),
    .Q_N(net797));
 sky130_fd_sc_hd__dfsbp_1 merge825 (.CLK(clknet_4_2_0_clk),
    .D(net302),
    .Q(net303),
    .Q_N(net799));
 sky130_fd_sc_hd__dfstp_1 merge826 (.CLK(clknet_4_3_0_clk),
    .D(net440),
    .SET_B(net738),
    .Q(net801));
 sky130_fd_sc_hd__dfstp_1 merge827 (.CLK(clknet_4_8_0_clk),
    .D(net757),
    .SET_B(net771),
    .Q(net802));
 sky130_fd_sc_hd__dfstp_1 merge828 (.CLK(clknet_4_2_0_clk),
    .D(net59),
    .Q(net60));
 sky130_fd_sc_hd__dlrbn_1 merge829 (.D(net566),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net577),
    .Q(net805),
    .Q_N(net804));
 sky130_fd_sc_hd__dlrbn_1 merge830 (.D(net316),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net325),
    .Q(net807),
    .Q_N(net806));
 sky130_fd_sc_hd__dlrbp_1 merge831 (.D(net540),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net739),
    .Q(net809),
    .Q_N(net808));
 sky130_fd_sc_hd__dlrbp_1 merge832 (.D(net488),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net492),
    .Q(net811),
    .Q_N(net810));
 sky130_fd_sc_hd__dlrtn_1 merge833 (.D(net653),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net654),
    .Q(net812));
 sky130_fd_sc_hd__dlrtn_1 merge834 (.GATE_N(clknet_4_10_0_clk),
    .RESET_B(net231),
    .Q(net232));
 sky130_fd_sc_hd__dlrtn_1 merge835 (.D(net429),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net431),
    .Q(net814));
 sky130_fd_sc_hd__dlrtp_1 merge836 (.D(net760),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net773),
    .Q(net815));
 sky130_fd_sc_hd__dlrtp_2 merge837 (.D(net258),
    .GATE(clknet_4_0_0_clk),
    .RESET_B(net260),
    .Q(net816));
 sky130_fd_sc_hd__dlrtp_1 merge838 (.D(net724),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net710),
    .Q(net817));
 sky130_fd_sc_hd__edfxbp_1 merge839 (.CLK(clknet_4_10_0_clk),
    .D(net98),
    .DE(net727),
    .Q(net819),
    .Q_N(net818));
 sky130_fd_sc_hd__edfxtp_1 merge840 (.CLK(clknet_4_7_0_clk),
    .D(net690),
    .DE(net708),
    .Q(net820));
 sky130_fd_sc_hd__sdlclkp_1 merge841 (.CLK(clknet_4_3_0_clk),
    .GATE(net562),
    .SCE(net544),
    .GCLK(net821));
 sky130_fd_sc_hd__sdlclkp_2 merge842 (.CLK(clknet_4_5_0_clk),
    .GATE(net633),
    .GCLK(net636));
 sky130_fd_sc_hd__sdlclkp_4 merge843 (.CLK(clknet_4_11_0_clk),
    .GATE(net335),
    .SCE(net342),
    .GCLK(net823));
 sky130_fd_sc_hd__dfrbp_1 merge844 (.CLK(clknet_4_7_0_clk),
    .D(net669),
    .RESET_B(net672),
    .Q(net825),
    .Q_N(net824));
 sky130_fd_sc_hd__dfrbp_1 merge845 (.CLK(clknet_4_12_0_clk),
    .D(net600),
    .RESET_B(net499),
    .Q(net826),
    .Q_N(net978));
 sky130_fd_sc_hd__and2_0 merge846 (.A(net661),
    .B(net588),
    .X(net827));
 sky130_fd_sc_hd__dfrtn_1 merge847 (.CLK_N(clknet_4_5_0_clk),
    .D(net673),
    .RESET_B(net682),
    .Q(net828));
 sky130_fd_sc_hd__dfrtp_1 merge848 (.CLK(clknet_4_10_0_clk),
    .D(net195),
    .RESET_B(net787),
    .Q(net829));
 sky130_fd_sc_hd__dfrtp_1 merge849 (.CLK(clknet_4_11_0_clk),
    .RESET_B(net793),
    .Q(net830));
 sky130_fd_sc_hd__dfrtp_2 merge850 (.CLK(clknet_4_4_0_clk),
    .D(net827),
    .RESET_B(net729),
    .Q(net831));
 sky130_fd_sc_hd__dfsbp_1 merge851 (.CLK(clknet_4_12_0_clk),
    .D(net607),
    .Q(net611),
    .Q_N(net832));
 sky130_fd_sc_hd__dfsbp_1 merge852 (.CLK(clknet_4_6_0_clk),
    .D(net579),
    .SET_B(net585),
    .Q(net835),
    .Q_N(net834));
 sky130_fd_sc_hd__dfstp_2 merge853 (.CLK(clknet_4_0_0_clk),
    .D(net764),
    .SET_B(net168),
    .Q(net836));
 sky130_fd_sc_hd__dfstp_1 merge854 (.CLK(clknet_4_8_0_clk),
    .D(net213),
    .SET_B(net745),
    .Q(net837));
 sky130_fd_sc_hd__dfstp_1 merge855 (.CLK(clknet_4_5_0_clk),
    .D(net674),
    .SET_B(net677),
    .Q(net838));
 sky130_fd_sc_hd__dlrbn_1 merge856 (.D(net713),
    .GATE_N(clknet_4_12_0_clk),
    .RESET_B(net476),
    .Q(net840),
    .Q_N(net839));
 sky130_fd_sc_hd__dlrbn_1 merge857 (.D(net493),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net498),
    .Q(net842),
    .Q_N(net841));
 sky130_fd_sc_hd__dlrbp_1 merge858 (.D(net281),
    .GATE(clknet_4_0_0_clk),
    .RESET_B(net282),
    .Q(net844),
    .Q_N(net843));
 sky130_fd_sc_hd__dlrbp_1 merge859 (.D(net582),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net496),
    .Q(net845),
    .Q_N(net967));
 sky130_fd_sc_hd__dlrtn_1 merge860 (.D(net786),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net765),
    .Q(net846));
 sky130_fd_sc_hd__dfxbp_2 s861 (.CLK(clknet_4_8_0_clk),
    .D(net57),
    .Q(net848),
    .Q_N(net847));
 sky130_fd_sc_hd__dfxbp_1 s862 (.CLK(clknet_4_8_0_clk),
    .D(net58),
    .Q(net850),
    .Q_N(net849));
 sky130_fd_sc_hd__dfxtp_1 s863 (.CLK(clknet_4_10_0_clk),
    .D(net70),
    .Q(net851));
 sky130_fd_sc_hd__dfxtp_1 s864 (.CLK(clknet_4_8_0_clk),
    .D(net82),
    .Q(net852));
 sky130_fd_sc_hd__dfxtp_1 s865 (.CLK(clknet_4_10_0_clk),
    .D(net100),
    .Q(net853));
 sky130_fd_sc_hd__dlclkp_1 s866 (.CLK(clknet_4_8_0_clk),
    .GATE(net190),
    .GCLK(net854));
 sky130_fd_sc_hd__dlclkp_2 s867 (.CLK(clknet_4_8_0_clk),
    .GATE(net192),
    .GCLK(net855));
 sky130_fd_sc_hd__dlclkp_4 s868 (.CLK(clknet_4_11_0_clk),
    .GATE(net215),
    .GCLK(net856));
 sky130_fd_sc_hd__dlxbn_2 s869 (.D(net293),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net858),
    .Q_N(net857));
 sky130_fd_sc_hd__dlxbn_1 s870 (.D(net296),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net860),
    .Q_N(net859));
 sky130_fd_sc_hd__dlxbp_1 s871 (.D(net298),
    .GATE(clknet_4_3_0_clk),
    .Q(net862),
    .Q_N(net861));
 sky130_fd_sc_hd__dlxtn_1 s872 (.D(net300),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net863));
 sky130_fd_sc_hd__dlxtn_1 s873 (.D(net317),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net864));
 sky130_fd_sc_hd__dlxtn_4 s874 (.D(net321),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net865));
 sky130_fd_sc_hd__dlxtp_1 s875 (.D(net326),
    .GATE(clknet_4_9_0_clk),
    .Q(net866));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s876 (.D(net343),
    .SLEEP_B(clknet_4_11_0_clk),
    .Q(net867));
 sky130_fd_sc_hd__dfxbp_1 s877 (.CLK(clknet_4_14_0_clk),
    .D(net345),
    .Q(net869),
    .Q_N(net868));
 sky130_fd_sc_hd__dfxbp_1 s878 (.CLK(clknet_4_11_0_clk),
    .D(net358),
    .Q(net871),
    .Q_N(net870));
 sky130_fd_sc_hd__dfxtp_1 s879 (.CLK(clknet_4_14_0_clk),
    .D(net369),
    .Q(net872));
 sky130_fd_sc_hd__dfxtp_1 s880 (.CLK(clknet_4_14_0_clk),
    .D(net372),
    .Q(net873));
 sky130_fd_sc_hd__dfxtp_1 s881 (.CLK(clknet_4_1_0_clk),
    .D(net412),
    .Q(net874));
 sky130_fd_sc_hd__dlclkp_1 s882 (.CLK(clknet_4_1_0_clk),
    .GATE(net413),
    .GCLK(net875));
 sky130_fd_sc_hd__dlclkp_2 s883 (.CLK(clknet_4_3_0_clk),
    .GATE(net435),
    .GCLK(net876));
 sky130_fd_sc_hd__dlclkp_4 s884 (.CLK(clknet_4_15_0_clk),
    .GATE(net456),
    .GCLK(net877));
 sky130_fd_sc_hd__dlxbn_1 s885 (.D(net473),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net879),
    .Q_N(net878));
 sky130_fd_sc_hd__dlxbn_1 s886 (.D(net482),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net881),
    .Q_N(net880));
 sky130_fd_sc_hd__dlxbp_1 s887 (.D(net490),
    .GATE(clknet_4_14_0_clk),
    .Q(net883),
    .Q_N(net882));
 sky130_fd_sc_hd__dlxtn_1 s888 (.D(net491),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net966));
 sky130_fd_sc_hd__dlxtn_1 s889 (.D(net495),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net970));
 sky130_fd_sc_hd__dlxtn_1 s890 (.D(net497),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net982));
 sky130_fd_sc_hd__dlxtp_1 s891 (.D(net516),
    .GATE(clknet_4_4_0_clk),
    .Q(net884));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s892 (.D(net523),
    .SLEEP_B(clknet_4_1_0_clk),
    .Q(net885));
 sky130_fd_sc_hd__dfxbp_1 s893 (.CLK(clknet_4_4_0_clk),
    .D(net539),
    .Q(net887),
    .Q_N(net886));
 sky130_fd_sc_hd__dfxbp_1 s894 (.CLK(clknet_4_4_0_clk),
    .D(net541),
    .Q(net889),
    .Q_N(net888));
 sky130_fd_sc_hd__dfxtp_2 s895 (.CLK(clknet_4_4_0_clk),
    .D(net542),
    .Q(net890));
 sky130_fd_sc_hd__dfxtp_1 s896 (.CLK(clknet_4_4_0_clk),
    .D(net549),
    .Q(net891));
 sky130_fd_sc_hd__dfxtp_1 s897 (.CLK(clknet_4_6_0_clk),
    .D(net561),
    .Q(net892));
 sky130_fd_sc_hd__dlclkp_1 s898 (.CLK(clknet_4_7_0_clk),
    .GATE(net584),
    .GCLK(net893));
 sky130_fd_sc_hd__dlclkp_2 s899 (.CLK(clknet_4_12_0_clk),
    .GATE(net604),
    .GCLK(net894));
 sky130_fd_sc_hd__dlclkp_4 s900 (.CLK(clknet_4_13_0_clk),
    .GATE(net610),
    .GCLK(net895));
 sky130_fd_sc_hd__dlxbn_1 s901 (.D(net612),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net896));
 sky130_fd_sc_hd__dlxbn_1 s902 (.D(net613),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net897));
 sky130_fd_sc_hd__dlxbp_1 s903 (.D(net614),
    .GATE(clknet_4_13_0_clk),
    .Q(net898));
 sky130_fd_sc_hd__dlxtn_1 s904 (.D(net657),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net899));
 sky130_fd_sc_hd__dlxtn_1 s905 (.D(net660),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net900));
 sky130_fd_sc_hd__dlxtn_1 s906 (.D(net662),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net901));
 sky130_fd_sc_hd__dlxtp_1 s907 (.D(net684),
    .GATE(clknet_4_7_0_clk),
    .Q(net902));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s908 (.D(net685),
    .SLEEP_B(clknet_4_7_0_clk),
    .Q(net903));
 sky130_fd_sc_hd__dfxbp_1 s909 (.CLK(clknet_4_7_0_clk),
    .D(net686),
    .Q(net905),
    .Q_N(net904));
 sky130_fd_sc_hd__dfxbp_1 s910 (.CLK(clknet_4_7_0_clk),
    .D(net689),
    .Q(net907),
    .Q_N(net906));
 sky130_fd_sc_hd__dfxtp_1 s911 (.CLK(clknet_4_7_0_clk),
    .D(net691),
    .Q(net908));
 sky130_fd_sc_hd__dfxtp_2 s912 (.CLK(clknet_4_7_0_clk),
    .D(net692),
    .Q(net909));
 sky130_fd_sc_hd__dfxtp_1 s913 (.CLK(clknet_4_7_0_clk),
    .D(net694),
    .Q(net910));
 sky130_fd_sc_hd__dlclkp_1 s914 (.CLK(clknet_4_7_0_clk),
    .GATE(net695),
    .GCLK(net911));
 sky130_fd_sc_hd__dlclkp_2 s915 (.CLK(clknet_4_7_0_clk),
    .GATE(net700),
    .GCLK(net912));
 sky130_fd_sc_hd__dlclkp_4 s916 (.CLK(clknet_4_7_0_clk),
    .GATE(net702),
    .GCLK(net913));
 sky130_fd_sc_hd__dlxbn_1 s917 (.D(net704),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net915),
    .Q_N(net914));
 sky130_fd_sc_hd__dlxbn_1 s918 (.D(net711),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net916));
 sky130_fd_sc_hd__dlxbp_1 s919 (.D(net714),
    .GATE(clknet_4_13_0_clk),
    .Q(net917));
 sky130_fd_sc_hd__dlxtn_1 s920 (.D(net715),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net918));
 sky130_fd_sc_hd__dlxtn_1 s921 (.D(net716),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net919));
 sky130_fd_sc_hd__dlxtn_1 s922 (.D(net718),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net920));
 sky130_fd_sc_hd__dlxtp_1 s923 (.D(net720),
    .GATE(clknet_4_13_0_clk),
    .Q(net921));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s924 (.D(net721),
    .SLEEP_B(clknet_4_13_0_clk),
    .Q(net922));
 sky130_fd_sc_hd__dfxbp_1 s925 (.CLK(clknet_4_13_0_clk),
    .D(net722),
    .Q(net923));
 sky130_fd_sc_hd__dfxbp_1 s926 (.CLK(clknet_4_0_0_clk),
    .D(net728),
    .Q(net925),
    .Q_N(net924));
 sky130_fd_sc_hd__dfxtp_1 s927 (.CLK(clknet_4_15_0_clk),
    .D(net733),
    .Q(net926));
 sky130_fd_sc_hd__dfxtp_1 s928 (.CLK(clknet_4_3_0_clk),
    .D(net736),
    .Q(net927));
 sky130_fd_sc_hd__dfxtp_1 s929 (.CLK(clknet_4_3_0_clk),
    .D(net740),
    .Q(net928));
 sky130_fd_sc_hd__dlclkp_1 s930 (.CLK(clknet_4_3_0_clk),
    .GATE(net746),
    .GCLK(net929));
 sky130_fd_sc_hd__dlclkp_2 s931 (.CLK(clknet_4_14_0_clk),
    .GATE(net747),
    .GCLK(net930));
 sky130_fd_sc_hd__dlclkp_4 s932 (.CLK(clknet_4_9_0_clk),
    .GATE(net761),
    .GCLK(net931));
 sky130_fd_sc_hd__dlxbn_1 s933 (.D(net767),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net933),
    .Q_N(net932));
 sky130_fd_sc_hd__dlxbn_1 s934 (.D(net770),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net935),
    .Q_N(net934));
 sky130_fd_sc_hd__dlxbp_1 s935 (.D(net772),
    .GATE(clknet_4_8_0_clk),
    .Q(net937),
    .Q_N(net936));
 sky130_fd_sc_hd__dlxtn_1 s936 (.D(net774),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net938));
 sky130_fd_sc_hd__dlxtn_1 s937 (.D(net775),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net939));
 sky130_fd_sc_hd__dlxtn_1 s938 (.D(net778),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net940));
 sky130_fd_sc_hd__dlxtp_1 s939 (.D(net779),
    .GATE(clknet_4_0_0_clk),
    .Q(net941));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s940 (.D(net781),
    .SLEEP_B(clknet_4_4_0_clk),
    .Q(net942));
 sky130_fd_sc_hd__dfxbp_1 s941 (.CLK(clknet_4_2_0_clk),
    .D(net782),
    .Q(net944),
    .Q_N(net943));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(in0),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(in1),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(in10),
    .X(net800));
 sky130_fd_sc_hd__buf_1 input4 (.A(in11),
    .X(net833));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(in12),
    .X(net945));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(in13),
    .X(net946));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(in14),
    .X(net947));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(in15),
    .X(net948));
 sky130_fd_sc_hd__buf_1 input9 (.A(in16),
    .X(net949));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(in17),
    .X(net950));
 sky130_fd_sc_hd__buf_1 input11 (.A(in18),
    .X(net951));
 sky130_fd_sc_hd__buf_1 input12 (.A(in19),
    .X(net952));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(in2),
    .X(net953));
 sky130_fd_sc_hd__buf_2 input14 (.A(in20),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(in21),
    .X(net955));
 sky130_fd_sc_hd__buf_2 input16 (.A(in22),
    .X(net956));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(in23),
    .X(net957));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(in24),
    .X(net958));
 sky130_fd_sc_hd__buf_1 input19 (.A(in3),
    .X(net959));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(in4),
    .X(net960));
 sky130_fd_sc_hd__buf_2 input21 (.A(in5),
    .X(net961));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(in6),
    .X(net962));
 sky130_fd_sc_hd__buf_4 input23 (.A(in7),
    .X(net963));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(in8),
    .X(net964));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(in9),
    .X(net965));
 sky130_fd_sc_hd__buf_2 output26 (.A(net966),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_4 output27 (.A(net967),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output28 (.A(net968),
    .X(out10));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(clknet_1_1__leaf_net969),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output30 (.A(net970),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output31 (.A(net971),
    .X(out13));
 sky130_fd_sc_hd__clkbuf_4 output32 (.A(net972),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output33 (.A(net973),
    .X(out15));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(clknet_1_1__leaf_net974),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output35 (.A(net975),
    .X(out17));
 sky130_fd_sc_hd__clkbuf_4 output36 (.A(net976),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output37 (.A(net977),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output38 (.A(net978),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output39 (.A(net979),
    .X(out20));
 sky130_fd_sc_hd__clkbuf_4 output40 (.A(net980),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output41 (.A(net981),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output42 (.A(net982),
    .X(out23));
 sky130_fd_sc_hd__clkbuf_1 output43 (.A(clknet_1_1__leaf_net983),
    .X(out24));
 sky130_fd_sc_hd__clkbuf_4 output44 (.A(net984),
    .X(out3));
 sky130_fd_sc_hd__clkbuf_1 output45 (.A(clknet_1_1__leaf_net985),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output46 (.A(net986),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output47 (.A(net987),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output48 (.A(net988),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_4 output49 (.A(net989),
    .X(out8));
 sky130_fd_sc_hd__clkbuf_4 output50 (.A(net990),
    .X(out9));
 sky130_fd_sc_hd__buf_4 fanout51 (.A(net256),
    .X(net991));
 sky130_fd_sc_hd__clkbuf_4 fanout52 (.A(net201),
    .X(net992));
 sky130_fd_sc_hd__buf_2 fanout53 (.A(net51),
    .X(net993));
 sky130_fd_sc_hd__clkbuf_4 fanout54 (.A(net280),
    .X(net994));
 sky130_fd_sc_hd__buf_2 fanout55 (.A(net996),
    .X(net995));
 sky130_fd_sc_hd__buf_2 fanout56 (.A(net997),
    .X(net996));
 sky130_fd_sc_hd__buf_8 fanout57 (.A(net161),
    .X(net997));
 sky130_fd_sc_hd__buf_12 fanout58 (.A(net145),
    .X(net998));
 sky130_fd_sc_hd__clkbuf_4 fanout59 (.A(net558),
    .X(net999));
 sky130_fd_sc_hd__clkbuf_2 fanout60 (.A(net558),
    .X(net1000));
 sky130_fd_sc_hd__buf_12 fanout61 (.A(net142),
    .X(net1001));
 sky130_fd_sc_hd__clkbuf_4 fanout62 (.A(net25),
    .X(net1002));
 sky130_fd_sc_hd__clkbuf_4 fanout63 (.A(net981),
    .X(net1003));
 sky130_fd_sc_hd__buf_2 fanout64 (.A(net642),
    .X(net1004));
 sky130_fd_sc_hd__clkbuf_4 fanout65 (.A(net626),
    .X(net1005));
 sky130_fd_sc_hd__buf_4 fanout66 (.A(net414),
    .X(net1006));
 sky130_fd_sc_hd__clkbuf_4 fanout67 (.A(net853),
    .X(net1007));
 sky130_fd_sc_hd__buf_2 fanout68 (.A(net355),
    .X(net1008));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net931 (.A(net931),
    .X(clknet_0_net931));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net931 (.A(clknet_0_net931),
    .X(clknet_1_0__leaf_net931));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net931 (.A(clknet_0_net931),
    .X(clknet_1_1__leaf_net931));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net329 (.A(net329),
    .X(clknet_0_net329));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net329 (.A(clknet_0_net329),
    .X(clknet_1_0__leaf_net329));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net329 (.A(clknet_0_net329),
    .X(clknet_1_1__leaf_net329));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net985 (.A(net985),
    .X(clknet_0_net985));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net985 (.A(clknet_0_net985),
    .X(clknet_1_0__leaf_net985));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net985 (.A(clknet_0_net985),
    .X(clknet_1_1__leaf_net985));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net361 (.A(net361),
    .X(clknet_0_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net361 (.A(clknet_0_net361),
    .X(clknet_1_0__leaf_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net361 (.A(net1036),
    .X(clknet_1_1__leaf_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net830 (.A(net830),
    .X(clknet_0_net830));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net830 (.A(clknet_0_net830),
    .X(clknet_1_0__leaf_net830));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net830 (.A(clknet_0_net830),
    .X(clknet_1_1__leaf_net830));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net338 (.A(net338),
    .X(clknet_0_net338));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net338 (.A(clknet_0_net338),
    .X(clknet_1_0__leaf_net338));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net338 (.A(clknet_0_net338),
    .X(clknet_1_1__leaf_net338));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net983 (.A(net983),
    .X(clknet_0_net983));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net983 (.A(clknet_0_net983),
    .X(clknet_1_0__leaf_net983));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net983 (.A(clknet_0_net983),
    .X(clknet_1_1__leaf_net983));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net292 (.A(net292),
    .X(clknet_0_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net292 (.A(clknet_0_net292),
    .X(clknet_1_0__leaf_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net292 (.A(clknet_0_net292),
    .X(clknet_1_1__leaf_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net427 (.A(net427),
    .X(clknet_0_net427));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net427 (.A(clknet_0_net427),
    .X(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net427 (.A(clknet_0_net427),
    .X(clknet_1_1__leaf_net427));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net929 (.A(net929),
    .X(clknet_0_net929));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net929 (.A(clknet_0_net929),
    .X(clknet_1_0__leaf_net929));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net929 (.A(clknet_0_net929),
    .X(clknet_1_1__leaf_net929));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net447 (.A(net447),
    .X(clknet_0_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net447 (.A(clknet_0_net447),
    .X(clknet_1_0__leaf_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net447 (.A(clknet_0_net447),
    .X(clknet_1_1__leaf_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net930 (.A(net930),
    .X(clknet_0_net930));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net930 (.A(clknet_0_net930),
    .X(clknet_1_0__leaf_net930));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net930 (.A(clknet_0_net930),
    .X(clknet_1_1__leaf_net930));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net451 (.A(net451),
    .X(clknet_0_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net451 (.A(clknet_0_net451),
    .X(clknet_1_0__leaf_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net451 (.A(clknet_0_net451),
    .X(clknet_1_1__leaf_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net481 (.A(net481),
    .X(clknet_0_net481));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net481 (.A(clknet_0_net481),
    .X(clknet_1_0__leaf_net481));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net481 (.A(clknet_0_net481),
    .X(clknet_1_1__leaf_net481));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net719 (.A(net719),
    .X(clknet_0_net719));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net719 (.A(clknet_0_net719),
    .X(clknet_1_0__leaf_net719));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net719 (.A(clknet_0_net719),
    .X(clknet_1_1__leaf_net719));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net593 (.A(net593),
    .X(clknet_0_net593));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net593 (.A(clknet_0_net593),
    .X(clknet_1_0__leaf_net593));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net593 (.A(clknet_0_net593),
    .X(clknet_1_1__leaf_net593));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net458 (.A(net458),
    .X(clknet_0_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net458 (.A(clknet_0_net458),
    .X(clknet_1_0__leaf_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net458 (.A(clknet_0_net458),
    .X(clknet_1_1__leaf_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net448 (.A(net448),
    .X(clknet_0_net448));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net448 (.A(clknet_0_net448),
    .X(clknet_1_0__leaf_net448));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net448 (.A(clknet_0_net448),
    .X(clknet_1_1__leaf_net448));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net877 (.A(net877),
    .X(clknet_0_net877));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net877 (.A(clknet_0_net877),
    .X(clknet_1_0__leaf_net877));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net877 (.A(clknet_0_net877),
    .X(clknet_1_1__leaf_net877));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net894 (.A(net894),
    .X(clknet_0_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net894 (.A(clknet_0_net894),
    .X(clknet_1_0__leaf_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net894 (.A(clknet_0_net894),
    .X(clknet_1_1__leaf_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net605 (.A(net605),
    .X(clknet_0_net605));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net605 (.A(clknet_0_net605),
    .X(clknet_1_0__leaf_net605));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net605 (.A(clknet_0_net605),
    .X(clknet_1_1__leaf_net605));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net567 (.A(net567),
    .X(clknet_0_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net567 (.A(clknet_0_net567),
    .X(clknet_1_0__leaf_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net567 (.A(clknet_0_net567),
    .X(clknet_1_1__leaf_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net609 (.A(net609),
    .X(clknet_0_net609));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net609 (.A(clknet_0_net609),
    .X(clknet_1_0__leaf_net609));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net609 (.A(clknet_0_net609),
    .X(clknet_1_1__leaf_net609));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net449 (.A(net449),
    .X(clknet_0_net449));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net449 (.A(clknet_0_net449),
    .X(clknet_1_0__leaf_net449));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net449 (.A(clknet_0_net449),
    .X(clknet_1_1__leaf_net449));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net457 (.A(net457),
    .X(clknet_0_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net457 (.A(clknet_0_net457),
    .X(clknet_1_0__leaf_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net457 (.A(clknet_0_net457),
    .X(clknet_1_1__leaf_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net911 (.A(net911),
    .X(clknet_0_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net911 (.A(clknet_0_net911),
    .X(clknet_1_0__leaf_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net911 (.A(clknet_0_net911),
    .X(clknet_1_1__leaf_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net707 (.A(net707),
    .X(clknet_0_net707));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net707 (.A(clknet_0_net707),
    .X(clknet_1_0__leaf_net707));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net707 (.A(clknet_0_net707),
    .X(clknet_1_1__leaf_net707));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net452 (.A(net452),
    .X(clknet_0_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net452 (.A(clknet_0_net452),
    .X(clknet_1_0__leaf_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net452 (.A(clknet_0_net452),
    .X(clknet_1_1__leaf_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net463 (.A(net463),
    .X(clknet_0_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net463 (.A(clknet_0_net463),
    .X(clknet_1_0__leaf_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net463 (.A(clknet_0_net463),
    .X(clknet_1_1__leaf_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net821 (.A(net821),
    .X(clknet_0_net821));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net821 (.A(clknet_0_net821),
    .X(clknet_1_0__leaf_net821));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net821 (.A(clknet_0_net821),
    .X(clknet_1_1__leaf_net821));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net546 (.A(net546),
    .X(clknet_0_net546));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net546 (.A(clknet_0_net546),
    .X(clknet_1_0__leaf_net546));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net546 (.A(clknet_0_net546),
    .X(clknet_1_1__leaf_net546));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net876 (.A(net876),
    .X(clknet_0_net876));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net876 (.A(clknet_0_net876),
    .X(clknet_1_0__leaf_net876));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net876 (.A(clknet_0_net876),
    .X(clknet_1_1__leaf_net876));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net436 (.A(net436),
    .X(clknet_0_net436));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net436 (.A(clknet_0_net436),
    .X(clknet_1_0__leaf_net436));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net436 (.A(clknet_0_net436),
    .X(clknet_1_1__leaf_net436));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net895 (.A(net895),
    .X(clknet_0_net895));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net895 (.A(clknet_0_net895),
    .X(clknet_1_0__leaf_net895));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net895 (.A(clknet_0_net895),
    .X(clknet_1_1__leaf_net895));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net913 (.A(net913),
    .X(clknet_0_net913));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net913 (.A(clknet_0_net913),
    .X(clknet_1_0__leaf_net913));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net913 (.A(clknet_0_net913),
    .X(clknet_1_1__leaf_net913));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net709 (.A(net709),
    .X(clknet_0_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net709 (.A(clknet_0_net709),
    .X(clknet_1_0__leaf_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net709 (.A(clknet_0_net709),
    .X(clknet_1_1__leaf_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net912 (.A(net912),
    .X(clknet_0_net912));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net912 (.A(clknet_0_net912),
    .X(clknet_1_0__leaf_net912));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net912 (.A(clknet_0_net912),
    .X(clknet_1_1__leaf_net912));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net893 (.A(net893),
    .X(clknet_0_net893));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net893 (.A(clknet_0_net893),
    .X(clknet_1_0__leaf_net893));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net893 (.A(clknet_0_net893),
    .X(clknet_1_1__leaf_net893));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net875 (.A(net875),
    .X(clknet_0_net875));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net875 (.A(clknet_0_net875),
    .X(clknet_1_0__leaf_net875));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net875 (.A(clknet_0_net875),
    .X(clknet_1_1__leaf_net875));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net420 (.A(net420),
    .X(clknet_0_net420));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net420 (.A(clknet_0_net420),
    .X(clknet_1_0__leaf_net420));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net420 (.A(clknet_0_net420),
    .X(clknet_1_1__leaf_net420));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net464 (.A(net464),
    .X(clknet_0_net464));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net464 (.A(clknet_0_net464),
    .X(clknet_1_0__leaf_net464));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net464 (.A(clknet_0_net464),
    .X(clknet_1_1__leaf_net464));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net424 (.A(net424),
    .X(clknet_0_net424));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net424 (.A(clknet_0_net424),
    .X(clknet_1_0__leaf_net424));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net424 (.A(clknet_0_net424),
    .X(clknet_1_1__leaf_net424));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net856 (.A(net856),
    .X(clknet_0_net856));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net856 (.A(clknet_0_net856),
    .X(clknet_1_0__leaf_net856));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net856 (.A(clknet_0_net856),
    .X(clknet_1_1__leaf_net856));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net353 (.A(net353),
    .X(clknet_0_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net353 (.A(clknet_0_net353),
    .X(clknet_1_0__leaf_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net353 (.A(clknet_0_net353),
    .X(clknet_1_1__leaf_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net221 (.A(net221),
    .X(clknet_0_net221));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net221 (.A(clknet_0_net221),
    .X(clknet_1_0__leaf_net221));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net221 (.A(clknet_0_net221),
    .X(clknet_1_1__leaf_net221));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net855 (.A(net855),
    .X(clknet_0_net855));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net855 (.A(clknet_0_net855),
    .X(clknet_1_0__leaf_net855));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net855 (.A(clknet_0_net855),
    .X(clknet_1_1__leaf_net855));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net823 (.A(net823),
    .X(clknet_0_net823));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net823 (.A(clknet_0_net823),
    .X(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net823 (.A(clknet_0_net823),
    .X(clknet_1_1__leaf_net823));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net346 (.A(net346),
    .X(clknet_0_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net346 (.A(clknet_0_net346),
    .X(clknet_1_0__leaf_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net346 (.A(clknet_0_net346),
    .X(clknet_1_1__leaf_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net974 (.A(net974),
    .X(clknet_0_net974));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net974 (.A(clknet_0_net974),
    .X(clknet_1_0__leaf_net974));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net974 (.A(clknet_0_net974),
    .X(clknet_1_1__leaf_net974));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net354 (.A(net354),
    .X(clknet_0_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net354 (.A(clknet_0_net354),
    .X(clknet_1_0__leaf_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net354 (.A(net1028),
    .X(clknet_1_1__leaf_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net854 (.A(net854),
    .X(clknet_0_net854));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net854 (.A(clknet_0_net854),
    .X(clknet_1_0__leaf_net854));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net854 (.A(clknet_0_net854),
    .X(clknet_1_1__leaf_net854));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net969 (.A(net969),
    .X(clknet_0_net969));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net969 (.A(clknet_0_net969),
    .X(clknet_1_0__leaf_net969));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net969 (.A(clknet_0_net969),
    .X(clknet_1_1__leaf_net969));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net315 (.A(net315),
    .X(clknet_0_net315));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net315 (.A(clknet_0_net315),
    .X(clknet_1_0__leaf_net315));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net315 (.A(clknet_0_net315),
    .X(clknet_1_1__leaf_net315));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net979),
    .X(net1009));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer2 (.A(net1009),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net979),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net160),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net1012),
    .X(net1013));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer6 (.A(net1013),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net1012),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net160),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net142),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net145),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net998),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net1019),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net1019),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net1019),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net1019),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net1001),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net1024),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net1025),
    .X(net1026));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer19 (.A(net1026),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(clknet_0_net354),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net237),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net237),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net17),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net1031),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net1031),
    .X(net1033));
 sky130_fd_sc_hd__clkbuf_1 clone26 (.A(net1035),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(net161),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(clknet_0_net361),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net852),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net794),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net872),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net834),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net938),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net804),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net859),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net791),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net873),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net909),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net99),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net842),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net814),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net1007),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net851),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net230),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net857),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net749),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net869),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net884),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net262),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net891),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net565),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net559),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net892),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net351),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net229),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net897),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net889),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net888),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net438),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net1004),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net675),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net925),
    .X(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_X (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_C_N (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S0 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_B (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_C1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_X (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_RESET_B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c39_C1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_X (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_C1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_D_N (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A0 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_S0 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_X (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_D (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_B (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_C1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A0 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_C1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_C (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_D_N (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_X (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_C1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_D (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A0 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_C1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_D_N (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_X (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_C (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_X (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_RESET_B (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_B (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_D_N (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A3 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_X (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_A0 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A0 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_C (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S0 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_SCE (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_B (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_C_N (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_X (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_C (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_X (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c47_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c39_X (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_C (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_S0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A3 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_SCD (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_X (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_C1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_X (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A3 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_X (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_B (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_RESET_B (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_X (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_C_N (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_RESET_B (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_A0 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_X (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A3 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_D (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_X (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_RESET_B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_C_N (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A0 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_X (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_D (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_X (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_A0 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_S0 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_C (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_X (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_A3 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A0 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_S0 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_D (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_X (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_SCD (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S0 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A3 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_C_N (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_D (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_S0 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_X (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_SCD (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_D1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A0 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_C_N (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_S1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A3 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_SCE (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_X (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_C_N (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_C (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_X (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_D (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_C1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A3 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_X (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_S0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_X (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_C (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_C1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_X (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_SCD (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_A3 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_D (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_D1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_SET_B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_SCD (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_D_N (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_SCD (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_X (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_RESET_B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_X (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_SCE (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_S1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_SCD (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_B (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_S0 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_X (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_S0 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_X (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold55_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A3 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_D1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_C_N (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A2 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_Q (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S0 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c53_B (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c49_X (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A0 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_A3 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_C1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A3 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_X (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_SCD (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S0 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_X (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S0 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_C_N (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_C (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_X (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A3 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c51_X (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_SCD (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_S0 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_D_N (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_X (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_C1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_S1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_X (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold49_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A0 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_D1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_C_N (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_C (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_X (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_S0 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_SET_B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S0 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A0 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_DE (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A3 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_C (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_X (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_D (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_RESET_B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_RESET_B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_X (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_C (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A3 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_D_N (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_C (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_X (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_C_N (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_S1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_C (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_C1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_X (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_RESET_B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c54_X (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_B1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_X (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_A2 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_A2 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_SCE (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_C (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A2 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_B (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_X (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A0 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A0 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_C (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_B1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_X (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_B1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_S0 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A0 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_C (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_X (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_S0 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_RESET_B (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_B (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_S1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A3 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_X (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_D (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_C (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_X (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_S1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c32_B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c28_X (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_B (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_S1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_S1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_C (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_SCE (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_C1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_X (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A0 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A3 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_B (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_D1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_C (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_X (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_SET_B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_S0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c60_C (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c57_X (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A0 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_X (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A0 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_X (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A3 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_B (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_D1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A3 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_X (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_C1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_C1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A0 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_B (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A3 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_B (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_X (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_X (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_A3 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_A (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_C1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_Q (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_S0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_X (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_S0 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_S0 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_B1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_SET_B (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_X (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_SCE (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_SCD (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_C (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_B (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S0 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_B (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_X (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_C_N (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_D (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_B (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_C (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_X (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_A2 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A2 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_X (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_X (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_SCE (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_B (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_B (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_X (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_B (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A3 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_B (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_C (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_X (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_C (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_X (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_D_N (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_B (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_C (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_B (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A3 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_X (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_A3 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_A3 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A3 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_RESET_B (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S1 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A3 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_SET_B (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_X (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_RESET_B (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_D_N (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_X (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_B (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_X (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_B (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A3 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_C (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_B (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A2 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_X (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_S1 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A2 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A1 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_C_N (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_SCD (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_B (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_X (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_B1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_C1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_SCD (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_Q_N (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold59_A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_Q (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_S0 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_SCE (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A2 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_X (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_C1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_D_N (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_X (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_D (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_S0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_SCE (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c35_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c30_X (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_C_N (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_A3 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_RESET_B (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A3 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_B (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_B (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_D (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_B (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_X (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_C_N (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_X (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S0 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A2 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_C (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A3 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S1 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_B (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_X (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_C1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A0 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_X (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_D_N (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_D (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_SCD (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A1 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_X (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S0 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A1 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_B (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_X (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_S1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_C_N (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_C (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_X (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A3 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_X (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_B (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_A0 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_SCD (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_SCD (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_B (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S0 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A3 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_X (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold52_A (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A0 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_Q (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net567_A (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_X (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S1 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_C1 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S1 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_D_N (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_Q_N (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_B1 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_Q (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c44_B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_A3 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_C1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c31_X (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_SCD (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A3 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_B (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_SCE (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_SCE (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_C (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_X (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_X (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout65_A (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S0 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_X (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_A2 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S0 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A1 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_C1 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A2 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_C (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_B1 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_B (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_X (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_A1 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S1 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A1 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_SET_B (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A3 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_B (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_X (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A0 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_SET_B (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_X (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_A (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A0 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_X (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A0 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A2 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_C1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_SCD (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_S0 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_C1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_B1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_X (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_C1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_X (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_RESET_B (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_X (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_B (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_Q (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_SET_B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_SCE (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_X (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A3 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_SCD (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_D_N (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A3 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_S1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_X (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_S1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_X (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_D1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A0 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_C1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_SCE (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_Q (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_RESET_B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_RESET_B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_X (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_X (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_Q (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_SCD (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_D1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_Q_N (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c39_B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_S0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c33_X (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_C (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_SCE (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A3 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_X (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_Q (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_D_N (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_SCE (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_C (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_C (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge850_Q (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A2 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_Q (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_SCD (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_Q_N (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_S0 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_B (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_s861_Q_N (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_B (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_D1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_S1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_D1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_S1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_s861_Q (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A2 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_C1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_D1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S0 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_B (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold45_A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_s869_Q_N (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A3 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_SCE (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_SCE (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S0 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_s869_Q (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S0 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_C1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_C_N (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_C1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_D1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_S0 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_S1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_s871_Q_N (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_S0 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_D1 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_D1 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_s871_Q (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_D_N (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_C (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_C (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_s874_Q (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A3 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_D1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_D1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_SCE (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_D_N (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_C (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_s881_Q (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_D1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_SET_B (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_B (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_Q (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_SET_B (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_SCE (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_Q (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_D1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_C (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_s908_Q (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S0 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S0 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S0 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_C1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold38_A (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_Q (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S0 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S1 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_B1 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A2 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S1 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S0 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S0 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_C1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A3 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_D1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_SCD (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_SCE (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_X (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_A3 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_X (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_RESET_B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_D_N (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_SET_B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_SET_B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_RESET_B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A3 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_X (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold39_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_C1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A3 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_X (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_B (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_C_N (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A0 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_RESET_B (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_B (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_B1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_A (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c51_B (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_D_N (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_SCD (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_C (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A2 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_RESET_B (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_C_N (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c30_B (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_A0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c46_A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_B (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_D_N (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_S1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c45_A (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_C_N (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A2 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_A1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c28_A (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_A1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_A (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_B (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_C_N (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_B (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c55_A (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_S0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_A3 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c27_B (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_B (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_C_N (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_SCE (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_B (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_S1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_A (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_C (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_SCD (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_C1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_C (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_B (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_output28_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_SCD (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_D (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_SCD (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_B1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_X (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_output32_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_A1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A2 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c61_C (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S0 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c58_X (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_B (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_output33_A (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_RESET_B (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_B (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_X (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_S0 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_B (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_B (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A3 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_X (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_output36_A (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_B (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_D_N (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_B1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_B1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_DE (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_S0 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_X (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_A (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_output41_A (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_A0 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_X (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_output44_A (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A2 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A3 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_C (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_X (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_output46_A (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_C1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_B (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_X (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_output48_A (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_SCE (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_B1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_A2 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_Q (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_output49_A (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_Q (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_output50_A (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_Q (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_X (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A3 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A3 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_D1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_B (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_S1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S0 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_D_N (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_X (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_B1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_S0 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_SCE (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_C_N (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_D1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_C1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A0 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_SCD (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A3 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_X (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_B (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_D_N (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_SCD (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_S1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_B (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_B (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_B (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_X (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_B (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_B (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A3 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_C (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A3 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A3 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_B (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A3 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout56_X (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_C (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_C (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_SET_B (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_S0 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_C_N (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout55_A (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout57_X (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_S0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_B1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_B (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout56_A (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_D1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer11_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_X (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_RESET_B (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_X (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_B (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_D_N (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_SET_B (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_C_N (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_DE (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_C1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer16_A (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_D1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_X (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_B1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_B (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_B (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_D_N (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_D_N (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_X (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_C (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S0 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A3 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c55_B (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c54_C (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c52_A (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_X (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_SCE (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_RESET_B (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_D_N (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold60_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_X (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_C1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_B1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_C1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A3 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_C1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_SCD (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_C_N (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_C (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout65_X (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A0 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S0 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A2 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_B1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_SCD (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_C_N (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_B (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_X (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A3 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_SCE (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_D_N (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_S0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_C (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold42_A (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout67_X (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_D1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_S1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_D1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_S1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_D1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_SCE (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_S1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_C_N (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s869_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s926_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s939_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge828_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s870_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s872_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s933_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s941_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s871_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s883_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s929_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge850_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s940_SLEEP_B (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge847_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s905_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s908_SLEEP_B (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s910_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s911_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge854_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s861_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s862_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s864_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s866_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s867_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s935_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s873_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s874_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s875_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s868_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_SLEEP_B (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s878_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s921_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s922_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s924_SLEEP_B (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s877_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s879_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s880_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_GATE (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge832_GATE (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_X (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_S1 (.DIODE(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_D_N (.DIODE(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S0 (.DIODE(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_S0 (.DIODE(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_DE (.DIODE(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A1 (.DIODE(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_A2 (.DIODE(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net427_X (.DIODE(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S1 (.DIODE(clknet_1_0__leaf_net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_D1 (.DIODE(clknet_1_0__leaf_net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_D1 (.DIODE(clknet_1_0__leaf_net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S1 (.DIODE(clknet_1_0__leaf_net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_D1 (.DIODE(clknet_1_0__leaf_net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net877_X (.DIODE(clknet_1_0__leaf_net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_B (.DIODE(clknet_1_0__leaf_net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_B (.DIODE(clknet_1_0__leaf_net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(clknet_1_0__leaf_net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net420_X (.DIODE(clknet_1_0__leaf_net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_SCD (.DIODE(clknet_1_1__leaf_net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(clknet_1_1__leaf_net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A1 (.DIODE(clknet_1_1__leaf_net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net420_X (.DIODE(clknet_1_1__leaf_net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_A (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_B (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_B (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_X (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_B (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_A (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A2 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer5_A (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_B1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer4_X (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer9_X (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_B (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer10_X (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer15_A (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer14_A (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_B (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer13_A (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_SCE (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer12_A (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer11_X (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone26_A (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer27_X (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_SET_B (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_S1 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold42_X (.DIODE(net1050));
 sky130_fd_sc_hd__and2_1 clone1 (.A(net946),
    .B(net955),
    .X(net1071));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
