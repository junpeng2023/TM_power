module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in62,
    in63,
    in64,
    in65,
    in66,
    in67,
    in68,
    in69,
    in7,
    in70,
    in71,
    in72,
    in73,
    in74,
    in75,
    in76,
    in77,
    in78,
    in79,
    in8,
    in80,
    in81,
    in82,
    in83,
    in84,
    in85,
    in86,
    in87,
    in88,
    in89,
    in9,
    in90,
    in91,
    in92,
    in93,
    in94,
    in95,
    in96,
    in97,
    in98,
    in99,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out62,
    out63,
    out64,
    out65,
    out66,
    out67,
    out68,
    out69,
    out7,
    out70,
    out71,
    out72,
    out73,
    out74,
    out75,
    out76,
    out77,
    out78,
    out79,
    out8,
    out80,
    out81,
    out82,
    out83,
    out84,
    out85,
    out86,
    out87,
    out88,
    out89,
    out9,
    out90,
    out91,
    out92,
    out93,
    out94,
    out95,
    out96,
    out97,
    out98,
    out99,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in62;
 input in63;
 input in64;
 input in65;
 input in66;
 input in67;
 input in68;
 input in69;
 input in7;
 input in70;
 input in71;
 input in72;
 input in73;
 input in74;
 input in75;
 input in76;
 input in77;
 input in78;
 input in79;
 input in8;
 input in80;
 input in81;
 input in82;
 input in83;
 input in84;
 input in85;
 input in86;
 input in87;
 input in88;
 input in89;
 input in9;
 input in90;
 input in91;
 input in92;
 input in93;
 input in94;
 input in95;
 input in96;
 input in97;
 input in98;
 input in99;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out62;
 output out63;
 output out64;
 output out65;
 output out66;
 output out67;
 output out68;
 output out69;
 output out7;
 output out70;
 output out71;
 output out72;
 output out73;
 output out74;
 output out75;
 output out76;
 output out77;
 output out78;
 output out79;
 output out8;
 output out80;
 output out81;
 output out82;
 output out83;
 output out84;
 output out85;
 output out86;
 output out87;
 output out88;
 output out89;
 output out9;
 output out90;
 output out91;
 output out92;
 output out93;
 output out94;
 output out95;
 output out96;
 output out97;
 output out98;
 output out99;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net412;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_0_net820;
 wire clknet_1_0__leaf_net820;
 wire clknet_1_1__leaf_net820;
 wire clknet_0_net529;
 wire clknet_1_0__leaf_net529;
 wire clknet_1_1__leaf_net529;
 wire clknet_0_net859;
 wire clknet_1_0__leaf_net859;
 wire clknet_1_1__leaf_net859;
 wire clknet_0_net523;
 wire clknet_1_0__leaf_net523;
 wire clknet_1_1__leaf_net523;
 wire clknet_0_net860;
 wire clknet_1_0__leaf_net860;
 wire clknet_1_1__leaf_net860;
 wire clknet_0_net539;
 wire clknet_1_0__leaf_net539;
 wire clknet_1_1__leaf_net539;
 wire clknet_0_net564;
 wire clknet_1_0__leaf_net564;
 wire clknet_1_1__leaf_net564;
 wire clknet_0_net681;
 wire clknet_1_0__leaf_net681;
 wire clknet_1_1__leaf_net681;
 wire clknet_0_net516;
 wire clknet_1_0__leaf_net516;
 wire clknet_1_1__leaf_net516;
 wire clknet_0_net992;
 wire clknet_1_0__leaf_net992;
 wire clknet_1_1__leaf_net992;
 wire clknet_0_net406;
 wire clknet_1_0__leaf_net406;
 wire clknet_1_1__leaf_net406;
 wire clknet_0_net651;
 wire clknet_1_0__leaf_net651;
 wire clknet_1_1__leaf_net651;
 wire clknet_0_net819;
 wire clknet_1_0__leaf_net819;
 wire clknet_1_1__leaf_net819;
 wire clknet_0_net391;
 wire clknet_1_0__leaf_net391;
 wire clknet_1_1__leaf_net391;
 wire clknet_0_net858;
 wire clknet_1_0__leaf_net858;
 wire clknet_1_1__leaf_net858;
 wire clknet_0_net818;
 wire clknet_1_0__leaf_net818;
 wire clknet_1_1__leaf_net818;
 wire clknet_0_net488;
 wire clknet_1_0__leaf_net488;
 wire clknet_1_1__leaf_net488;
 wire clknet_0_net394;
 wire clknet_1_0__leaf_net394;
 wire clknet_1_1__leaf_net394;
 wire clknet_0_net393;
 wire clknet_1_0__leaf_net393;
 wire clknet_1_1__leaf_net393;
 wire clknet_0_net839;
 wire clknet_1_0__leaf_net839;
 wire clknet_1_1__leaf_net839;
 wire clknet_0_net464;
 wire clknet_1_0__leaf_net464;
 wire clknet_1_1__leaf_net464;
 wire clknet_0_net462;
 wire clknet_1_0__leaf_net462;
 wire clknet_1_1__leaf_net462;
 wire clknet_0_net970;
 wire clknet_1_0__leaf_net970;
 wire clknet_1_1__leaf_net970;
 wire clknet_0_net390;
 wire clknet_1_0__leaf_net390;
 wire clknet_1_1__leaf_net390;
 wire clknet_0_net389;
 wire clknet_1_0__leaf_net389;
 wire clknet_1_1__leaf_net389;
 wire clknet_0_net387;
 wire clknet_1_0__leaf_net387;
 wire clknet_1_1__leaf_net387;
 wire clknet_0_net802;
 wire clknet_1_0__leaf_net802;
 wire clknet_1_1__leaf_net802;
 wire clknet_0_net1000;
 wire clknet_1_0__leaf_net1000;
 wire clknet_1_1__leaf_net1000;
 wire clknet_0_net341;
 wire clknet_1_0__leaf_net341;
 wire clknet_1_1__leaf_net341;
 wire clknet_0_net332;
 wire clknet_1_0__leaf_net332;
 wire clknet_1_1__leaf_net332;
 wire clknet_0_net331;
 wire clknet_1_0__leaf_net331;
 wire clknet_1_1__leaf_net331;
 wire clknet_0_net340;
 wire clknet_1_0__leaf_net340;
 wire clknet_1_1__leaf_net340;
 wire clknet_0_net801;
 wire clknet_1_0__leaf_net801;
 wire clknet_1_1__leaf_net801;
 wire clknet_0_net431;
 wire clknet_1_0__leaf_net431;
 wire clknet_1_1__leaf_net431;
 wire clknet_0_net365;
 wire clknet_1_0__leaf_net365;
 wire clknet_1_1__leaf_net365;
 wire clknet_0_net460;
 wire clknet_1_0__leaf_net460;
 wire clknet_1_1__leaf_net460;
 wire clknet_0_net458;
 wire clknet_1_0__leaf_net458;
 wire clknet_1_1__leaf_net458;
 wire clknet_0_net324;
 wire clknet_1_0__leaf_net324;
 wire clknet_1_1__leaf_net324;
 wire clknet_0_net328;
 wire clknet_1_0__leaf_net328;
 wire clknet_1_1__leaf_net328;
 wire clknet_0_net800;
 wire clknet_1_0__leaf_net800;
 wire clknet_1_1__leaf_net800;
 wire clknet_0_net425;
 wire clknet_1_0__leaf_net425;
 wire clknet_1_1__leaf_net425;
 wire clknet_0_net439;
 wire clknet_1_0__leaf_net439;
 wire clknet_1_1__leaf_net439;
 wire clknet_0_net838;
 wire clknet_1_0__leaf_net838;
 wire clknet_1_1__leaf_net838;
 wire clknet_0_net999;
 wire clknet_1_0__leaf_net999;
 wire clknet_1_1__leaf_net999;
 wire clknet_0_net493;
 wire clknet_1_0__leaf_net493;
 wire clknet_1_1__leaf_net493;
 wire clknet_0_net784;
 wire clknet_1_0__leaf_net784;
 wire clknet_1_1__leaf_net784;
 wire clknet_0_net783;
 wire clknet_1_0__leaf_net783;
 wire clknet_1_1__leaf_net783;
 wire clknet_0_net396;
 wire clknet_1_0__leaf_net396;
 wire clknet_1_1__leaf_net396;
 wire clknet_0_net969;
 wire clknet_1_0__leaf_net969;
 wire clknet_1_1__leaf_net969;
 wire clknet_0_net301;
 wire clknet_1_0__leaf_net301;
 wire clknet_1_1__leaf_net301;
 wire clknet_0_net782;
 wire clknet_1_0__leaf_net782;
 wire clknet_1_1__leaf_net782;
 wire clknet_0_net361;
 wire clknet_1_0__leaf_net361;
 wire clknet_1_1__leaf_net361;
 wire clknet_0_net976;
 wire clknet_1_0__leaf_net976;
 wire clknet_1_1__leaf_net976;
 wire clknet_0_net290;
 wire clknet_1_0__leaf_net290;
 wire clknet_1_1__leaf_net290;
 wire clknet_0_net287;
 wire clknet_1_0__leaf_net287;
 wire clknet_1_1__leaf_net287;
 wire clknet_0_net296;
 wire clknet_1_0__leaf_net296;
 wire clknet_1_1__leaf_net296;
 wire clknet_0_net291;
 wire clknet_1_0__leaf_net291;
 wire clknet_1_1__leaf_net291;
 wire clknet_0_net279;
 wire clknet_1_0__leaf_net279;
 wire clknet_1_1__leaf_net279;
 wire clknet_0_net766;
 wire clknet_1_0__leaf_net766;
 wire clknet_1_1__leaf_net766;
 wire clknet_0_net637;
 wire clknet_1_0__leaf_net637;
 wire clknet_1_1__leaf_net637;
 wire clknet_0_net990;
 wire clknet_1_0__leaf_net990;
 wire clknet_1_1__leaf_net990;
 wire clknet_0_net840;
 wire clknet_1_0__leaf_net840;
 wire clknet_1_1__leaf_net840;
 wire clknet_0_net456;
 wire clknet_1_0__leaf_net456;
 wire clknet_1_1__leaf_net456;
 wire clknet_0_net223;
 wire clknet_1_0__leaf_net223;
 wire clknet_1_1__leaf_net223;
 wire clknet_0_net1022;
 wire clknet_1_0__leaf_net1022;
 wire clknet_1_1__leaf_net1022;
 wire clknet_0_net325;
 wire clknet_1_0__leaf_net325;
 wire clknet_1_1__leaf_net325;
 wire clknet_0_net765;
 wire clknet_1_0__leaf_net765;
 wire clknet_1_1__leaf_net765;
 wire clknet_0_net346;
 wire clknet_1_0__leaf_net346;
 wire clknet_1_1__leaf_net346;
 wire clknet_0_net996;
 wire clknet_1_0__leaf_net996;
 wire clknet_1_1__leaf_net996;
 wire clknet_0_net435;
 wire clknet_1_0__leaf_net435;
 wire clknet_1_1__leaf_net435;
 wire clknet_0_net214;
 wire clknet_1_0__leaf_net214;
 wire clknet_1_1__leaf_net214;
 wire clknet_0_net202;
 wire clknet_1_0__leaf_net202;
 wire clknet_1_1__leaf_net202;
 wire clknet_0_net764;
 wire clknet_1_0__leaf_net764;
 wire clknet_1_1__leaf_net764;
 wire clknet_0_net232;
 wire clknet_1_0__leaf_net232;
 wire clknet_1_1__leaf_net232;
 wire clknet_0_net233;
 wire clknet_1_0__leaf_net233;
 wire clknet_1_1__leaf_net233;
 wire clknet_0_net745;
 wire clknet_1_0__leaf_net745;
 wire clknet_1_1__leaf_net745;
 wire clknet_0_net257;
 wire clknet_1_0__leaf_net257;
 wire clknet_1_1__leaf_net257;
 wire clknet_0_net255;
 wire clknet_1_0__leaf_net255;
 wire clknet_1_1__leaf_net255;
 wire clknet_0_net261;
 wire clknet_1_0__leaf_net261;
 wire clknet_1_1__leaf_net261;
 wire clknet_0_net256;
 wire clknet_1_0__leaf_net256;
 wire clknet_1_1__leaf_net256;
 wire clknet_0_net269;
 wire clknet_1_0__leaf_net269;
 wire clknet_1_1__leaf_net269;
 wire clknet_0_net744;
 wire clknet_1_0__leaf_net744;
 wire clknet_1_1__leaf_net744;
 wire clknet_0_net430;
 wire clknet_1_0__leaf_net430;
 wire clknet_1_1__leaf_net430;
 wire clknet_0_net398;
 wire clknet_1_0__leaf_net398;
 wire clknet_1_1__leaf_net398;
 wire clknet_0_net400;
 wire clknet_1_0__leaf_net400;
 wire clknet_1_1__leaf_net400;
 wire clknet_0_net1002;
 wire clknet_1_0__leaf_net1002;
 wire clknet_1_1__leaf_net1002;
 wire clknet_0_net211;
 wire clknet_1_0__leaf_net211;
 wire clknet_1_1__leaf_net211;
 wire clknet_0_net215;
 wire clknet_1_0__leaf_net215;
 wire clknet_1_1__leaf_net215;
 wire clknet_0_net743;
 wire clknet_1_0__leaf_net743;
 wire clknet_1_1__leaf_net743;
 wire clknet_0_net503;
 wire clknet_1_0__leaf_net503;
 wire clknet_1_1__leaf_net503;
 wire clknet_0_net513;
 wire clknet_1_0__leaf_net513;
 wire clknet_1_1__leaf_net513;
 wire clknet_0_net525;
 wire clknet_1_0__leaf_net525;
 wire clknet_1_1__leaf_net525;
 wire clknet_0_net519;
 wire clknet_1_0__leaf_net519;
 wire clknet_1_1__leaf_net519;
 wire clknet_0_net506;
 wire clknet_1_0__leaf_net506;
 wire clknet_1_1__leaf_net506;
 wire clknet_0_net505;
 wire clknet_1_0__leaf_net505;
 wire clknet_1_1__leaf_net505;
 wire clknet_0_net504;
 wire clknet_1_0__leaf_net504;
 wire clknet_1_1__leaf_net504;
 wire clknet_0_net185;
 wire clknet_1_0__leaf_net185;
 wire clknet_1_1__leaf_net185;
 wire clknet_0_net193;
 wire clknet_1_0__leaf_net193;
 wire clknet_1_1__leaf_net193;
 wire clknet_0_net191;
 wire clknet_1_0__leaf_net191;
 wire clknet_1_1__leaf_net191;
 wire clknet_0_net189;
 wire clknet_1_0__leaf_net189;
 wire clknet_1_1__leaf_net189;
 wire clknet_0_net197;
 wire clknet_1_0__leaf_net197;
 wire clknet_1_1__leaf_net197;
 wire clknet_0_net164;
 wire clknet_1_0__leaf_net164;
 wire clknet_1_1__leaf_net164;
 wire clknet_0_net726;
 wire clknet_1_0__leaf_net726;
 wire clknet_1_1__leaf_net726;
 wire clknet_0_net725;
 wire clknet_1_0__leaf_net725;
 wire clknet_1_1__leaf_net725;
 wire clknet_0_net112;
 wire clknet_1_0__leaf_net112;
 wire clknet_1_1__leaf_net112;
 wire clknet_0_net102;
 wire clknet_1_0__leaf_net102;
 wire clknet_1_1__leaf_net102;
 wire clknet_0_net987;
 wire clknet_1_0__leaf_net987;
 wire clknet_1_1__leaf_net987;
 wire clknet_0_net117;
 wire clknet_1_0__leaf_net117;
 wire clknet_1_1__leaf_net117;
 wire clknet_0_net113;
 wire clknet_1_0__leaf_net113;
 wire clknet_1_1__leaf_net113;
 wire clknet_0_net100;
 wire clknet_1_0__leaf_net100;
 wire clknet_1_1__leaf_net100;
 wire clknet_0_net104;
 wire clknet_1_0__leaf_net104;
 wire clknet_1_1__leaf_net104;
 wire clknet_0_net206;
 wire clknet_1_0__leaf_net206;
 wire clknet_1_1__leaf_net206;
 wire clknet_0_net103;
 wire clknet_1_0__leaf_net103;
 wire clknet_1_1__leaf_net103;
 wire clknet_0_net724;
 wire clknet_1_0__leaf_net724;
 wire clknet_1_1__leaf_net724;
 wire clknet_0_net705;
 wire clknet_1_0__leaf_net705;
 wire clknet_1_1__leaf_net705;
 wire clknet_0_net181;
 wire clknet_1_0__leaf_net181;
 wire clknet_1_1__leaf_net181;
 wire clknet_0_net404;
 wire clknet_1_0__leaf_net404;
 wire clknet_1_1__leaf_net404;
 wire clknet_0_net183;
 wire clknet_1_0__leaf_net183;
 wire clknet_1_1__leaf_net183;
 wire clknet_0_net88;
 wire clknet_1_0__leaf_net88;
 wire clknet_1_1__leaf_net88;
 wire clknet_0_net635;
 wire clknet_1_0__leaf_net635;
 wire clknet_1_1__leaf_net635;
 wire clknet_0_net1003;
 wire clknet_1_0__leaf_net1003;
 wire clknet_1_1__leaf_net1003;
 wire clknet_0_net82;
 wire clknet_1_0__leaf_net82;
 wire clknet_1_1__leaf_net82;
 wire clknet_0_net83;
 wire clknet_1_0__leaf_net83;
 wire clknet_1_1__leaf_net83;
 wire clknet_0_net979;
 wire clknet_1_0__leaf_net979;
 wire clknet_1_1__leaf_net979;
 wire clknet_0_net704;
 wire clknet_1_0__leaf_net704;
 wire clknet_1_1__leaf_net704;
 wire clknet_0_net217;
 wire clknet_1_0__leaf_net217;
 wire clknet_1_1__leaf_net217;
 wire clknet_0_net241;
 wire clknet_1_0__leaf_net241;
 wire clknet_1_1__leaf_net241;
 wire clknet_0_net225;
 wire clknet_1_0__leaf_net225;
 wire clknet_1_1__leaf_net225;
 wire clknet_0_net703;
 wire clknet_1_0__leaf_net703;
 wire clknet_1_1__leaf_net703;
 wire clknet_0_net277;
 wire clknet_1_0__leaf_net277;
 wire clknet_1_1__leaf_net277;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;

 sky130_fd_sc_hd__mux4_2 c100 (.A0(net958),
    .A1(net960),
    .A2(net955),
    .A3(net1126),
    .S0(net965),
    .S1(net936),
    .X(net0));
 sky130_fd_sc_hd__mux4_1 c101 (.A0(net952),
    .A1(net965),
    .A2(net960),
    .A3(net958),
    .S0(net959),
    .S1(net936),
    .X(net1));
 sky130_fd_sc_hd__mux4_2 c102 (.A0(net1122),
    .A1(net959),
    .A2(net960),
    .A3(net932),
    .S0(net950),
    .S1(net965),
    .X(net1021));
 sky130_fd_sc_hd__mux4_2 c103 (.A0(net960),
    .A1(net952),
    .A2(net959),
    .A3(net965),
    .S0(net961),
    .S1(net918),
    .X(net1042));
 sky130_fd_sc_hd__mux4_1 c104 (.A0(net1),
    .A1(net939),
    .A2(net955),
    .A3(net965),
    .S0(net951),
    .S1(net942),
    .X(net2));
 sky130_fd_sc_hd__mux4_2 c105 (.A0(net965),
    .A1(net960),
    .A2(net2),
    .A3(net959),
    .S0(net961),
    .S1(net1104),
    .X(net3));
 sky130_fd_sc_hd__mux4_1 c106 (.A0(net956),
    .A1(net961),
    .A2(net3),
    .A3(net939),
    .S0(net916),
    .S1(net1125),
    .X(net4));
 sky130_fd_sc_hd__mux4_2 c107 (.A0(net959),
    .A1(net939),
    .A2(net958),
    .A3(net934),
    .S0(net965),
    .S1(net1023),
    .X(net1008));
 sky130_fd_sc_hd__mux4_1 c108 (.A0(net2),
    .A1(net884),
    .A2(net966),
    .A3(net961),
    .S0(net938),
    .S1(net1008),
    .X(net5));
 sky130_fd_sc_hd__mux4_1 c109 (.A0(net967),
    .A1(net939),
    .A2(net5),
    .A3(net3),
    .S0(net887),
    .S1(net1008),
    .X(net6));
 sky130_fd_sc_hd__mux4_1 c110 (.A0(net1),
    .A1(net958),
    .A2(net921),
    .A3(net1021),
    .S0(net918),
    .S1(net1113),
    .X(net7));
 sky130_fd_sc_hd__a41o_1 c111 (.A1(net893),
    .A2(net934),
    .A3(net922),
    .A4(net7),
    .B1(net1095),
    .X(net8));
 sky130_fd_sc_hd__a41o_1 c112 (.A1(net918),
    .A2(net945),
    .A3(net887),
    .A4(net1),
    .B1(net1113),
    .X(net9));
 sky130_fd_sc_hd__a41o_2 c113 (.A1(net956),
    .A2(net936),
    .A3(net950),
    .A4(net912),
    .B1(net922),
    .X(net1019));
 sky130_fd_sc_hd__a41o_1 c114 (.A1(net9),
    .A2(net2),
    .A3(net912),
    .A4(net1096),
    .B1(net950),
    .X(net1032));
 sky130_fd_sc_hd__mux4_1 c115 (.A0(net958),
    .A1(net934),
    .A2(net1019),
    .A3(net961),
    .S0(net1113),
    .S1(net1096),
    .X(net1041));
 sky130_fd_sc_hd__a41o_1 c116 (.A1(net887),
    .A2(net8),
    .A3(net1042),
    .A4(net1041),
    .B1(net890),
    .X(net10));
 sky130_fd_sc_hd__mux4_1 c117 (.A0(net947),
    .A1(net963),
    .A2(net9),
    .A3(net1098),
    .S0(net1032),
    .S1(net921),
    .X(net11));
 sky130_fd_sc_hd__mux4_2 c118 (.A0(net936),
    .A1(net918),
    .A2(net1041),
    .A3(net1113),
    .S0(net9),
    .S1(net1031),
    .X(net12));
 sky130_fd_sc_hd__sdfbbn_1 c119 (.CLK_N(clknet_leaf_36_clk),
    .D(net1113),
    .RESET_B(net12),
    .SCD(net934),
    .SCE(net1107),
    .SET_B(net921),
    .Q(net14),
    .Q_N(net13));
 sky130_fd_sc_hd__a41o_1 c120 (.A1(net887),
    .A2(net1019),
    .A3(net1096),
    .A4(net921),
    .B1(net936),
    .X(net1044));
 sky130_fd_sc_hd__a41o_1 c121 (.A1(net950),
    .A2(net14),
    .A3(net904),
    .A4(net947),
    .B1(net964),
    .X(net1043));
 sky130_fd_sc_hd__a41o_1 c122 (.A1(net926),
    .A2(net915),
    .A3(net1044),
    .A4(net912),
    .B1(net1113),
    .X(net1034));
 sky130_fd_sc_hd__a41o_1 c123 (.A1(net7),
    .A2(net12),
    .A3(net1034),
    .A4(net13),
    .B1(net1044),
    .X(net15));
 sky130_fd_sc_hd__mux4_2 c124 (.A0(net1096),
    .A1(net887),
    .A2(net13),
    .A3(net921),
    .S0(net962),
    .S1(net1113),
    .X(net1026));
 sky130_fd_sc_hd__mux4_2 c125 (.A0(net963),
    .A1(net965),
    .A2(net912),
    .A3(net945),
    .S0(net950),
    .S1(net887),
    .X(net1017));
 sky130_fd_sc_hd__mux4_1 c126 (.A0(net14),
    .A1(net920),
    .A2(net918),
    .A3(net942),
    .S0(net1032),
    .S1(net1169),
    .X(net16));
 sky130_fd_sc_hd__mux4_2 c127 (.A0(net912),
    .A1(net1034),
    .A2(net1017),
    .A3(net950),
    .S0(net963),
    .S1(net1045),
    .X(net17));
 sky130_fd_sc_hd__a41o_1 c128 (.A1(net1019),
    .A2(net1034),
    .A3(net956),
    .A4(net1045),
    .B1(net1166),
    .X(net18));
 sky130_fd_sc_hd__a41o_1 c129 (.A1(net945),
    .A2(net1019),
    .A3(net1017),
    .A4(net13),
    .B1(net922),
    .X(net19));
 sky130_fd_sc_hd__mux4_1 c130 (.A0(net19),
    .A1(net947),
    .A2(net12),
    .A3(net1151),
    .S0(net1047),
    .S1(net1045),
    .X(net20));
 sky130_fd_sc_hd__mux4_1 c131 (.A0(net12),
    .A1(net1017),
    .A2(net964),
    .A3(net1008),
    .S0(net1026),
    .S1(net1149),
    .X(net21));
 sky130_fd_sc_hd__a41o_4 c132 (.A1(net1099),
    .A2(net1125),
    .A3(net1108),
    .A4(net1095),
    .B1(net1111),
    .X(net22));
 sky130_fd_sc_hd__a41o_2 c133 (.A1(net22),
    .A2(net1093),
    .A3(net1124),
    .A4(net1094),
    .B1(net1122),
    .X(net23));
 sky130_fd_sc_hd__a31o_2 c134 (.A1(net1124),
    .A2(net873),
    .A3(net1093),
    .B1(net1112),
    .X(net1039));
 sky130_fd_sc_hd__a41o_4 c135 (.A1(net873),
    .A2(net1095),
    .A3(net1092),
    .A4(net1125),
    .B1(net1098),
    .X(net24));
 sky130_fd_sc_hd__a41o_2 c136 (.A1(net24),
    .A2(net1074),
    .A3(net1107),
    .A4(net1111),
    .B1(net1117),
    .X(net25));
 sky130_fd_sc_hd__a31o_2 c137 (.A1(net1100),
    .A2(net22),
    .A3(net1102),
    .B1(net1111),
    .X(net26));
 sky130_fd_sc_hd__a41o_2 c138 (.A1(net1094),
    .A2(net1124),
    .A3(net1104),
    .A4(net24),
    .B1(net1074),
    .X(net968));
 sky130_fd_sc_hd__a41o_2 c139 (.A1(net24),
    .A2(net1095),
    .A3(net1106),
    .A4(net1074),
    .B1(net1073),
    .X(net27));
 sky130_fd_sc_hd__sdfbbn_2 c140 (.CLK_N(clknet_leaf_48_clk),
    .D(net1099),
    .RESET_B(net1111),
    .SCD(net1058),
    .SCE(net1060),
    .SET_B(net25),
    .Q(net29),
    .Q_N(net28));
 sky130_fd_sc_hd__a41o_1 c141 (.A1(net1073),
    .A2(net1104),
    .A3(net1058),
    .A4(net1111),
    .B1(net1090),
    .X(net30));
 sky130_fd_sc_hd__mux4_1 c142 (.A0(net870),
    .A1(net1094),
    .A2(net1060),
    .A3(net24),
    .S0(net1090),
    .S1(net611),
    .X(net31));
 sky130_fd_sc_hd__a41o_1 c143 (.A1(net870),
    .A2(net25),
    .A3(net1060),
    .A4(net1091),
    .B1(net1148),
    .X(net32));
 sky130_fd_sc_hd__mux4_1 c144 (.A0(net1058),
    .A1(net1060),
    .A2(net1111),
    .A3(net1090),
    .S0(net610),
    .S1(net697),
    .X(net33));
 sky130_fd_sc_hd__mux4_1 c145 (.A0(net1060),
    .A1(net1093),
    .A2(net1058),
    .A3(net1127),
    .S0(net1124),
    .S1(net699),
    .X(net34));
 sky130_fd_sc_hd__sdfbbp_1 c146 (.CLK(clknet_leaf_49_clk),
    .D(net25),
    .RESET_B(net1094),
    .SCD(net1090),
    .SCE(net698),
    .SET_B(net1144),
    .Q(net36),
    .Q_N(net35));
 sky130_fd_sc_hd__mux4_2 c147 (.A0(net24),
    .A1(net1124),
    .A2(net1074),
    .A3(net1111),
    .S0(net1090),
    .S1(net610),
    .X(net37));
 sky130_fd_sc_hd__sdfbbn_2 c148 (.CLK_N(clknet_leaf_49_clk),
    .D(net1057),
    .RESET_B(net1090),
    .SCD(net611),
    .SCE(net697),
    .SET_B(net698),
    .Q(net974),
    .Q_N(net38));
 sky130_fd_sc_hd__sdfbbn_2 c149 (.CLK_N(clknet_leaf_1_clk),
    .D(net1058),
    .RESET_B(net1091),
    .SCD(net974),
    .SCE(net611),
    .SET_B(net696),
    .Q(net40),
    .Q_N(net39));
 sky130_fd_sc_hd__mux4_2 c150 (.A0(net36),
    .A1(net870),
    .A2(net873),
    .A3(net1074),
    .S0(net38),
    .S1(net696),
    .X(net41));
 sky130_fd_sc_hd__sdfbbp_1 c151 (.CLK(clknet_leaf_49_clk),
    .D(net24),
    .RESET_B(net1057),
    .SCD(net39),
    .SCE(net1090),
    .SET_B(net1144),
    .Q(net983),
    .Q_N(net42));
 sky130_fd_sc_hd__mux4_1 c152 (.A0(net1095),
    .A1(net1056),
    .A2(net42),
    .A3(net1091),
    .S0(net1074),
    .S1(net39),
    .X(net43));
 sky130_fd_sc_hd__mux4_1 c153 (.A0(net983),
    .A1(net25),
    .A2(net1057),
    .A3(net611),
    .S0(net699),
    .S1(net1082),
    .X(net44));
 sky130_fd_sc_hd__a41o_2 c154 (.A1(net895),
    .A2(net1117),
    .A3(net1118),
    .A4(net1098),
    .B1(net1112),
    .X(net45));
 sky130_fd_sc_hd__mux4_2 c155 (.A0(net1124),
    .A1(net45),
    .A2(net896),
    .A3(net1120),
    .S0(net1118),
    .S1(net895),
    .X(net46));
 sky130_fd_sc_hd__sdfbbn_2 c156 (.CLK_N(clknet_leaf_44_clk),
    .D(net25),
    .RESET_B(net1095),
    .SCD(net46),
    .SCE(net38),
    .SET_B(net1073),
    .Q(net48),
    .Q_N(net47));
 sky130_fd_sc_hd__mux4_2 c157 (.A0(net1074),
    .A1(net888),
    .A2(net889),
    .A3(net1120),
    .S0(net890),
    .S1(net1118),
    .X(net49));
 sky130_fd_sc_hd__a41o_1 c158 (.A1(net45),
    .A2(net47),
    .A3(net38),
    .A4(net901),
    .B1(net611),
    .X(net50));
 sky130_fd_sc_hd__a41o_1 c159 (.A1(net896),
    .A2(net1093),
    .A3(net1071),
    .A4(net1095),
    .B1(net49),
    .X(net51));
 sky130_fd_sc_hd__sdfbbn_2 c160 (.CLK_N(clknet_leaf_46_clk),
    .D(net1125),
    .RESET_B(net1095),
    .SCD(net49),
    .SCE(net1071),
    .SET_B(net47),
    .Q(net1016),
    .Q_N(net52));
 sky130_fd_sc_hd__a41o_2 c161 (.A1(net1016),
    .A2(net45),
    .A3(net1071),
    .A4(net47),
    .B1(net598),
    .X(net53));
 sky130_fd_sc_hd__sdfbbp_1 c162 (.CLK(clknet_leaf_47_clk),
    .D(net1102),
    .RESET_B(net896),
    .SCD(net1100),
    .SCE(net49),
    .SET_B(net45),
    .Q(net1028),
    .Q_N(net54));
 sky130_fd_sc_hd__mux4_2 c163 (.A0(net873),
    .A1(net1016),
    .A2(net1109),
    .A3(net889),
    .S0(net1071),
    .S1(net47),
    .X(net55));
 sky130_fd_sc_hd__mux4_1 c164 (.A0(net1054),
    .A1(net901),
    .A2(net1120),
    .A3(net39),
    .S0(net1122),
    .S1(net895),
    .X(net56));
 sky130_fd_sc_hd__mux4_1 c165 (.A0(net1055),
    .A1(net1028),
    .A2(net1054),
    .A3(net870),
    .S0(net35),
    .S1(net1104),
    .X(net57));
 sky130_fd_sc_hd__sdfbbn_2 c166 (.CLK_N(clknet_leaf_7_clk),
    .D(net873),
    .RESET_B(net905),
    .SCD(net1093),
    .SCE(net1055),
    .SET_B(clknet_1_1__leaf_net704),
    .Q(net59),
    .Q_N(net58));
 sky130_fd_sc_hd__a41o_1 c167 (.A1(net59),
    .A2(net888),
    .A3(net1016),
    .A4(net1071),
    .B1(net46),
    .X(net60));
 sky130_fd_sc_hd__mux4_1 c168 (.A0(net1100),
    .A1(net25),
    .A2(net1054),
    .A3(net54),
    .S0(net60),
    .S1(clknet_1_0__leaf_net703),
    .X(net61));
 sky130_fd_sc_hd__mux4_1 c169 (.A0(net1071),
    .A1(net1028),
    .A2(net45),
    .A3(net889),
    .S0(net1100),
    .S1(clknet_1_0__leaf_net705),
    .X(net979));
 sky130_fd_sc_hd__mux4_1 c170 (.A0(net60),
    .A1(net1125),
    .A2(net896),
    .A3(net883),
    .S0(net903),
    .S1(net888),
    .X(net62));
 sky130_fd_sc_hd__mux4_1 c171 (.A0(net897),
    .A1(net1016),
    .A2(net1071),
    .A3(net1054),
    .S0(clknet_1_0__leaf_net703),
    .S1(net707),
    .X(net63));
 sky130_fd_sc_hd__mux4_1 c172 (.A0(net60),
    .A1(net46),
    .A2(net1055),
    .A3(net1085),
    .S0(clknet_1_0__leaf_net705),
    .S1(net706),
    .X(net64));
 sky130_fd_sc_hd__mux4_2 c173 (.A0(net889),
    .A1(net1107),
    .A2(net22),
    .A3(net1016),
    .S0(net598),
    .S1(net629),
    .X(net65));
 sky130_fd_sc_hd__a41o_1 c174 (.A1(net60),
    .A2(net1120),
    .A3(net1085),
    .B1(net706),
    .X(net66));
 sky130_fd_sc_hd__mux4_1 c175 (.A0(net1125),
    .A1(net1070),
    .A2(net60),
    .A3(net629),
    .S0(net1082),
    .S1(net707),
    .X(net67));
 sky130_fd_sc_hd__mux4_1 c176 (.A0(net928),
    .A1(net923),
    .A2(net917),
    .A3(net25),
    .S0(net1099),
    .S1(net1122),
    .X(net68));
 sky130_fd_sc_hd__mux4_1 c177 (.A0(net25),
    .A1(net897),
    .A2(net54),
    .A3(net1118),
    .S0(net42),
    .S1(net1070),
    .X(net69));
 sky130_fd_sc_hd__mux4_2 c178 (.A0(net919),
    .A1(net911),
    .A2(net1109),
    .A3(net908),
    .S0(net926),
    .S1(net920),
    .X(net70));
 sky130_fd_sc_hd__mux4_1 c179 (.A0(net1107),
    .A1(net917),
    .A2(net1056),
    .A3(net925),
    .S0(net1099),
    .S1(net710),
    .X(net71));
 sky130_fd_sc_hd__a41o_1 c180 (.A1(net1120),
    .A2(net929),
    .A3(net907),
    .A4(net926),
    .B1(net1127),
    .X(net72));
 sky130_fd_sc_hd__a41o_4 c181 (.A1(net901),
    .A2(net72),
    .A3(net898),
    .A4(net42),
    .B1(net712),
    .X(net73));
 sky130_fd_sc_hd__a41o_2 c182 (.A1(net1117),
    .A2(net925),
    .A3(net930),
    .A4(net910),
    .B1(net1099),
    .X(net74));
 sky130_fd_sc_hd__mux4_2 c183 (.A0(net1122),
    .A1(net928),
    .A2(net929),
    .A3(net917),
    .S0(net911),
    .S1(net919),
    .X(net986));
 sky130_fd_sc_hd__mux4_1 c184 (.A0(net888),
    .A1(net73),
    .A2(net1016),
    .A3(net72),
    .S0(net49),
    .S1(net713),
    .X(net75));
 sky130_fd_sc_hd__a41o_1 c185 (.A1(net72),
    .A2(net70),
    .A3(net1109),
    .A4(net712),
    .B1(net714),
    .X(net76));
 sky130_fd_sc_hd__mux4_2 c186 (.A0(net910),
    .A1(net48),
    .A2(net889),
    .A3(net38),
    .S0(net710),
    .S1(net713),
    .X(net77));
 sky130_fd_sc_hd__mux4_2 c187 (.A0(net889),
    .A1(net70),
    .A2(net915),
    .A3(net1126),
    .S0(net47),
    .S1(net713),
    .X(net78));
 sky130_fd_sc_hd__mux4_1 c188 (.A0(net60),
    .A1(net919),
    .A2(net78),
    .A3(net901),
    .S0(net713),
    .S1(net714),
    .X(net79));
 sky130_fd_sc_hd__mux4_2 c189 (.A0(net76),
    .A1(net909),
    .A2(net70),
    .A3(net1099),
    .S0(net78),
    .S1(net714),
    .X(net80));
 sky130_fd_sc_hd__mux4_1 c190 (.A0(net74),
    .A1(net80),
    .A2(net70),
    .A3(net1127),
    .S0(net612),
    .S1(net714),
    .X(net81));
 sky130_fd_sc_hd__mux4_1 c191 (.A0(net986),
    .A1(net1110),
    .A2(net919),
    .A3(net58),
    .S0(net1085),
    .S1(clknet_1_0__leaf_net635),
    .X(net82));
 sky130_fd_sc_hd__mux4_1 c192 (.A0(net78),
    .A1(net1091),
    .A2(clknet_1_0__leaf_net82),
    .A3(net919),
    .S0(net612),
    .S1(net707),
    .X(net83));
 sky130_fd_sc_hd__mux4_1 c193 (.A0(net926),
    .A1(clknet_1_0__leaf_net82),
    .A2(clknet_1_0__leaf_net83),
    .A3(net925),
    .S0(net930),
    .S1(net612),
    .X(net84));
 sky130_fd_sc_hd__mux4_1 c194 (.A0(net910),
    .A1(net901),
    .A2(clknet_1_0__leaf_net83),
    .A3(net80),
    .S0(clknet_1_0__leaf_net705),
    .S1(net715),
    .X(net85));
 sky130_fd_sc_hd__mux4_1 c195 (.A0(clknet_1_0__leaf_net83),
    .A1(net1091),
    .A2(net908),
    .A3(net74),
    .S0(clknet_1_0__leaf_net635),
    .S1(net715),
    .X(net86));
 sky130_fd_sc_hd__mux4_1 c196 (.A0(net927),
    .A1(clknet_1_0__leaf_net635),
    .A2(net712),
    .A3(net714),
    .S0(net715),
    .S1(net716),
    .X(net1003));
 sky130_fd_sc_hd__a41o_1 c197 (.A1(net80),
    .A2(net897),
    .A3(net1125),
    .B1(clknet_1_0__leaf_net635),
    .X(net87));
 sky130_fd_sc_hd__mux4_1 c198 (.A0(net933),
    .A1(net1110),
    .A2(net76),
    .A3(net1113),
    .S0(clknet_1_1__leaf_net703),
    .S1(clknet_1_0__leaf_net705),
    .X(net88));
 sky130_fd_sc_hd__mux4_1 c199 (.A0(net1104),
    .A1(net934),
    .A2(net1054),
    .A3(net1070),
    .S0(net1082),
    .S1(net714),
    .X(net89));
 sky130_fd_sc_hd__mux4_1 c200 (.A0(net80),
    .A1(net52),
    .A2(net953),
    .A3(net597),
    .S0(net697),
    .S1(net712),
    .X(net90));
 sky130_fd_sc_hd__mux4_1 c201 (.A0(net923),
    .A1(net936),
    .A2(clknet_1_0__leaf_net88),
    .A3(net598),
    .S0(net629),
    .S1(net696),
    .X(net91));
 sky130_fd_sc_hd__mux4_1 c202 (.A0(net916),
    .A1(clknet_1_0__leaf_net82),
    .A2(clknet_1_0__leaf_net88),
    .A3(net47),
    .S0(net923),
    .S1(net997),
    .X(net92));
 sky130_fd_sc_hd__mux4_1 c203 (.A0(net1123),
    .A1(net74),
    .A2(net941),
    .A3(clknet_1_1__leaf_net88),
    .S0(net1122),
    .S1(net1107),
    .X(net93));
 sky130_fd_sc_hd__mux4_1 c204 (.A0(net943),
    .A1(net931),
    .A2(net884),
    .A3(net916),
    .S0(clknet_1_0__leaf_net88),
    .S1(net720),
    .X(net94));
 sky130_fd_sc_hd__mux4_1 c205 (.A0(clknet_1_0__leaf_net88),
    .A1(net940),
    .A2(net1070),
    .A3(net1109),
    .S0(net1072),
    .S1(net722),
    .X(net95));
 sky130_fd_sc_hd__mux4_1 c206 (.A0(net933),
    .A1(net1110),
    .A2(net943),
    .A3(clknet_1_0__leaf_net88),
    .S0(net722),
    .S1(clknet_1_0__leaf_net724),
    .X(net96));
 sky130_fd_sc_hd__mux4_1 c207 (.A0(clknet_1_1__leaf_net82),
    .A1(clknet_1_0__leaf_net88),
    .A2(net718),
    .A3(net719),
    .S0(net722),
    .S1(net723),
    .X(net97));
 sky130_fd_sc_hd__mux4_1 c208 (.A0(net888),
    .A1(clknet_1_0__leaf_net88),
    .A2(net937),
    .A3(net1113),
    .S0(clknet_1_0__leaf_net724),
    .S1(clknet_1_0__leaf_net726),
    .X(net98));
 sky130_fd_sc_hd__mux4_1 c209 (.A0(net1127),
    .A1(clknet_1_0__leaf_net88),
    .A2(clknet_1_0__leaf_net635),
    .A3(net713),
    .S0(clknet_1_0__leaf_net725),
    .S1(clknet_1_1__leaf_net726),
    .X(net99));
 sky130_fd_sc_hd__mux4_2 c210 (.A0(net938),
    .A1(net612),
    .A2(net713),
    .A3(net720),
    .S0(net723),
    .S1(clknet_1_0__leaf_net725),
    .X(net100));
 sky130_fd_sc_hd__mux4_1 c211 (.A0(net936),
    .A1(net36),
    .A2(clknet_1_1__leaf_net88),
    .A3(net76),
    .S0(net906),
    .S1(clknet_1_0__leaf_net635),
    .X(net101));
 sky130_fd_sc_hd__mux4_1 c212 (.A0(clknet_1_0__leaf_net100),
    .A1(net909),
    .A2(net954),
    .A3(net696),
    .S0(clknet_1_1__leaf_net725),
    .S1(net729),
    .X(net102));
 sky130_fd_sc_hd__mux4_1 c213 (.A0(net944),
    .A1(net46),
    .A2(clknet_1_0__leaf_net100),
    .A3(net915),
    .S0(net719),
    .S1(net721),
    .X(net103));
 sky130_fd_sc_hd__mux4_1 c214 (.A0(net927),
    .A1(net890),
    .A2(clknet_1_0__leaf_net100),
    .A3(net997),
    .S0(net717),
    .S1(clknet_1_1__leaf_net724),
    .X(net104));
 sky130_fd_sc_hd__mux4_1 c215 (.A0(net953),
    .A1(clknet_1_0__leaf_net103),
    .A2(net70),
    .A3(clknet_1_0__leaf_net100),
    .S0(net944),
    .S1(net612),
    .X(net105));
 sky130_fd_sc_hd__mux4_1 c216 (.A0(net930),
    .A1(clknet_1_0__leaf_net104),
    .A2(clknet_1_0__leaf_net88),
    .A3(net884),
    .S0(net612),
    .S1(clknet_1_0__leaf_net726),
    .X(net106));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(clknet_1_0__leaf_net100),
    .A1(net1060),
    .A2(net884),
    .A3(clknet_1_0__leaf_net103),
    .S0(net728),
    .S1(net732),
    .X(net107));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(net70),
    .A1(clknet_1_0__leaf_net104),
    .A2(clknet_1_0__leaf_net88),
    .A3(clknet_1_0__leaf_net100),
    .S0(clknet_1_0__leaf_net726),
    .S1(net732),
    .X(net108));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net936),
    .A1(net22),
    .A2(net1092),
    .A3(clknet_1_0__leaf_net88),
    .S0(net732),
    .S1(net1077),
    .X(net109));
 sky130_fd_sc_hd__mux4_1 c220 (.A0(net1113),
    .A1(net73),
    .A2(net942),
    .A3(clknet_1_0__leaf_net83),
    .S0(clknet_1_0__leaf_net88),
    .S1(net730),
    .X(net110));
 sky130_fd_sc_hd__mux4_1 c221 (.A0(net1092),
    .A1(net3),
    .A2(net1070),
    .A3(net931),
    .S0(net1126),
    .S1(net598),
    .X(net111));
 sky130_fd_sc_hd__mux4_2 c222 (.A0(net932),
    .A1(net955),
    .A2(net1092),
    .A3(net960),
    .S0(net1023),
    .S1(net729),
    .X(net1035));
 sky130_fd_sc_hd__mux4_1 c223 (.A0(net0),
    .A1(net1102),
    .A2(net960),
    .A3(net1125),
    .S0(net35),
    .S1(clknet_1_1__leaf_net725),
    .X(net112));
 sky130_fd_sc_hd__mux4_1 c224 (.A0(net1089),
    .A1(net934),
    .A2(clknet_1_0__leaf_net102),
    .A3(net1125),
    .S0(net1081),
    .S1(clknet_1_1__leaf_net703),
    .X(net113));
 sky130_fd_sc_hd__mux4_1 c225 (.A0(net884),
    .A1(net1122),
    .A2(clknet_1_0__leaf_net113),
    .A3(net931),
    .S0(net1042),
    .S1(net927),
    .X(net114));
 sky130_fd_sc_hd__mux4_1 c226 (.A0(net77),
    .A1(net1008),
    .A2(net893),
    .A3(clknet_1_1__leaf_net88),
    .S0(net1081),
    .S1(clknet_1_1__leaf_net705),
    .X(net115));
 sky130_fd_sc_hd__mux4_1 c227 (.A0(net955),
    .A1(net1061),
    .A2(net52),
    .A3(net1107),
    .S0(net922),
    .S1(net734),
    .X(net116));
 sky130_fd_sc_hd__mux4_1 c228 (.A0(net951),
    .A1(net986),
    .A2(net1121),
    .A3(net38),
    .S0(net1023),
    .S1(net734),
    .X(net1025));
 sky130_fd_sc_hd__mux4_1 c229 (.A0(clknet_1_0__leaf_net102),
    .A1(net1109),
    .A2(net951),
    .A3(net52),
    .S0(net734),
    .S1(net737),
    .X(net117));
 sky130_fd_sc_hd__mux4_1 c230 (.A0(clknet_1_1__leaf_net102),
    .A1(net922),
    .A2(net52),
    .A3(net77),
    .S0(net1004),
    .S1(net1077),
    .X(net987));
 sky130_fd_sc_hd__mux4_1 c231 (.A0(net931),
    .A1(net881),
    .A2(clknet_1_0__leaf_net987),
    .A3(net723),
    .S0(net1077),
    .S1(net737),
    .X(net118));
 sky130_fd_sc_hd__mux4_1 c232 (.A0(clknet_1_0__leaf_net117),
    .A1(net73),
    .A2(clknet_1_0__leaf_net112),
    .A3(net1114),
    .S0(net710),
    .S1(net735),
    .X(net119));
 sky130_fd_sc_hd__mux4_1 c233 (.A0(net1125),
    .A1(clknet_1_0__leaf_net117),
    .A2(clknet_1_0__leaf_net112),
    .A3(net1042),
    .S0(clknet_1_0__leaf_net987),
    .S1(net735),
    .X(net120));
 sky130_fd_sc_hd__mux4_1 c234 (.A0(net0),
    .A1(net942),
    .A2(net1114),
    .A3(clknet_1_0__leaf_net88),
    .S0(net738),
    .S1(net740),
    .X(net121));
 sky130_fd_sc_hd__mux4_1 c235 (.A0(net939),
    .A1(clknet_1_1__leaf_net117),
    .A2(clknet_1_0__leaf_net987),
    .A3(clknet_1_1__leaf_net102),
    .S0(net619),
    .S1(net740),
    .X(net122));
 sky130_fd_sc_hd__mux4_1 c236 (.A0(net938),
    .A1(clknet_1_0__leaf_net88),
    .A2(net1021),
    .A3(net1004),
    .S0(net712),
    .S1(net735),
    .X(net123));
 sky130_fd_sc_hd__mux4_1 c237 (.A0(net78),
    .A1(net1121),
    .A2(clknet_1_0__leaf_net987),
    .A3(net1081),
    .S0(net732),
    .S1(net741),
    .X(net124));
 sky130_fd_sc_hd__mux4_2 c238 (.A0(net939),
    .A1(net38),
    .A2(net712),
    .A3(net730),
    .S0(net739),
    .S1(net740),
    .X(net1038));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net1038),
    .A1(net967),
    .A2(net878),
    .A3(net633),
    .S0(net716),
    .S1(net723),
    .X(net125));
 sky130_fd_sc_hd__mux4_1 c240 (.A0(net942),
    .A1(net1118),
    .A2(net125),
    .A3(net633),
    .S0(net683),
    .S1(net735),
    .X(net1027));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(net5),
    .A1(net1027),
    .A2(net1038),
    .A3(net1025),
    .S0(net125),
    .S1(net1161),
    .X(net126));
 sky130_fd_sc_hd__mux4_1 c256 (.A0(net8),
    .A1(net1043),
    .A2(net1099),
    .A3(net893),
    .S0(net1023),
    .S1(net738),
    .X(net127));
 sky130_fd_sc_hd__mux4_1 c257 (.A0(net942),
    .A1(net14),
    .A2(net8),
    .A3(net1038),
    .S0(net1019),
    .S1(net934),
    .X(net128));
 sky130_fd_sc_hd__mux4_1 c258 (.A0(net967),
    .A1(clknet_1_0__leaf_net987),
    .A2(net1023),
    .A3(net683),
    .S0(net1036),
    .S1(net742),
    .X(net129));
 sky130_fd_sc_hd__mux4_1 c259 (.A0(net14),
    .A1(net1035),
    .A2(net1026),
    .A3(net1038),
    .S0(net1092),
    .S1(net742),
    .X(net1037));
 sky130_fd_sc_hd__mux4_1 c260 (.A0(net125),
    .A1(net893),
    .A2(net942),
    .A3(net962),
    .S0(net1042),
    .S1(net742),
    .X(net1024));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(net926),
    .A1(net1043),
    .A2(clknet_1_0__leaf_net1003),
    .A3(net1037),
    .S0(clknet_1_0__leaf_net987),
    .S1(net742),
    .X(net130));
 sky130_fd_sc_hd__mux4_1 c262 (.A0(clknet_1_1__leaf_net117),
    .A1(net1037),
    .A2(net961),
    .A3(net1018),
    .S0(net711),
    .S1(net742),
    .X(net131));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net967),
    .A1(net903),
    .A2(net1046),
    .A3(net1018),
    .S0(net1031),
    .S1(net711),
    .X(net1048));
 sky130_fd_sc_hd__a41o_2 c264 (.A1(net1095),
    .A2(net1073),
    .A3(net24),
    .A4(net610),
    .B1(net698),
    .X(net132));
 sky130_fd_sc_hd__sdfbbn_2 c265 (.CLK_N(clknet_leaf_1_clk),
    .D(net1106),
    .RESET_B(net22),
    .SCD(net1092),
    .SCE(net1111),
    .SET_B(net1056),
    .Q(net1006),
    .Q_N(net133));
 sky130_fd_sc_hd__a41o_1 c266 (.A1(net1117),
    .A2(net133),
    .A3(net1121),
    .A4(net1090),
    .B1(net696),
    .X(net134));
 sky130_fd_sc_hd__sdfbbp_1 c267 (.CLK(clknet_leaf_50_clk),
    .D(net1108),
    .RESET_B(net1066),
    .SCD(net1122),
    .SCE(net132),
    .SET_B(net1144),
    .Q(net136),
    .Q_N(net135));
 sky130_fd_sc_hd__sdfbbn_2 c268 (.CLK_N(clknet_leaf_1_clk),
    .D(net1094),
    .RESET_B(net132),
    .SCD(net1123),
    .SCE(net1067),
    .SET_B(net1056),
    .Q(net138),
    .Q_N(net137));
 sky130_fd_sc_hd__a41o_1 c269 (.A1(net132),
    .A2(net133),
    .A3(net1066),
    .A4(net1094),
    .B1(net1148),
    .X(net139));
 sky130_fd_sc_hd__sdfbbn_2 c270 (.CLK_N(clknet_leaf_0_clk),
    .D(net138),
    .RESET_B(net1066),
    .SCD(net132),
    .SCE(net1100),
    .SET_B(net700),
    .Q(net141),
    .Q_N(net140));
 sky130_fd_sc_hd__sdfbbp_1 c271 (.CLK(clknet_leaf_0_clk),
    .D(net132),
    .RESET_B(net1074),
    .SCD(net1066),
    .SCE(net1167),
    .SET_B(net1080),
    .Q(net143),
    .Q_N(net142));
 sky130_fd_sc_hd__a41o_1 c272 (.A1(net1104),
    .A2(net1087),
    .A3(net1066),
    .A4(net611),
    .B1(net617),
    .X(net144));
 sky130_fd_sc_hd__a41o_1 c273 (.A1(net144),
    .A2(net136),
    .A3(net1067),
    .A4(net1086),
    .B1(net38),
    .X(net145));
 sky130_fd_sc_hd__mux4_2 c274 (.A0(net1122),
    .A1(net141),
    .A2(net1091),
    .A3(net1121),
    .S0(net1086),
    .S1(net1066),
    .X(net146));
 sky130_fd_sc_hd__sdfbbn_2 c275 (.CLK_N(clknet_leaf_0_clk),
    .D(net145),
    .RESET_B(net873),
    .SCD(net1086),
    .SCE(net140),
    .SET_B(net1067),
    .Q(net148),
    .Q_N(net147));
 sky130_fd_sc_hd__mux4_2 c276 (.A0(net1126),
    .A1(net144),
    .A2(net140),
    .A3(net1104),
    .S0(net1086),
    .S1(net1067),
    .X(net149));
 sky130_fd_sc_hd__a41o_1 c277 (.A1(net1006),
    .A2(net1087),
    .A3(net1067),
    .A4(net1053),
    .B1(net617),
    .X(net150));
 sky130_fd_sc_hd__sdfbbn_2 c278 (.CLK_N(clknet_leaf_0_clk),
    .D(net149),
    .RESET_B(net1087),
    .SCD(net1095),
    .SCE(net145),
    .SET_B(net1066),
    .Q(net152),
    .Q_N(net151));
 sky130_fd_sc_hd__a41o_2 c279 (.A1(net1123),
    .A2(net148),
    .A3(net1066),
    .A4(net22),
    .B1(net1086),
    .X(net153));
 sky130_fd_sc_hd__a41o_1 c280 (.A1(net870),
    .A2(net1087),
    .A3(net1053),
    .A4(net140),
    .B1(net1066),
    .X(net154));
 sky130_fd_sc_hd__mux4_1 c281 (.A0(net150),
    .A1(net151),
    .A2(net1086),
    .A3(net1050),
    .S0(net1111),
    .S1(net617),
    .X(net155));
 sky130_fd_sc_hd__mux4_1 c282 (.A0(net145),
    .A1(net1050),
    .A2(net1086),
    .A3(net1066),
    .S0(net610),
    .S1(clknet_1_0__leaf_net743),
    .X(net156));
 sky130_fd_sc_hd__mux4_1 c283 (.A0(net152),
    .A1(net144),
    .A2(net1050),
    .A3(net1086),
    .S0(net617),
    .S1(clknet_1_0__leaf_net743),
    .X(net157));
 sky130_fd_sc_hd__mux4_1 c284 (.A0(net141),
    .A1(net149),
    .A2(net1087),
    .A3(net1050),
    .S0(net1053),
    .S1(clknet_1_0__leaf_net743),
    .X(net158));
 sky130_fd_sc_hd__mux4_1 c285 (.A0(net149),
    .A1(net1050),
    .A2(net151),
    .A3(net870),
    .S0(clknet_1_0__leaf_net744),
    .S1(clknet_1_0__leaf_net745),
    .X(net159));
 sky130_fd_sc_hd__mux4_1 c286 (.A0(net1107),
    .A1(net1108),
    .A2(net1054),
    .A3(net1093),
    .S0(net629),
    .S1(clknet_1_0__leaf_net703),
    .X(net160));
 sky130_fd_sc_hd__sdfbbp_1 c287 (.CLK(clknet_leaf_5_clk),
    .D(net906),
    .RESET_B(net1052),
    .SCD(net153),
    .SCE(net629),
    .SET_B(clknet_1_0__leaf_net703),
    .Q(net162),
    .Q_N(net161));
 sky130_fd_sc_hd__a41o_4 c288 (.A1(net45),
    .A2(net1087),
    .A3(net35),
    .A4(net58),
    .B1(net1080),
    .X(net163));
 sky130_fd_sc_hd__a41o_1 c289 (.A1(net883),
    .A2(net163),
    .A3(net1070),
    .A4(net895),
    .B1(clknet_1_0__leaf_net743),
    .X(net164));
 sky130_fd_sc_hd__mux4_2 c290 (.A0(net1109),
    .A1(net1124),
    .A2(net1112),
    .A3(net893),
    .S0(net883),
    .S1(net1080),
    .X(net165));
 sky130_fd_sc_hd__sdfbbn_2 c291 (.CLK_N(clknet_leaf_2_clk),
    .D(net890),
    .RESET_B(net1164),
    .SCD(net135),
    .SCE(net1056),
    .SET_B(net1142),
    .Q(net167),
    .Q_N(net166));
 sky130_fd_sc_hd__mux4_1 c292 (.A0(net167),
    .A1(net904),
    .A2(net163),
    .A3(net1124),
    .S0(net132),
    .S1(net629),
    .X(net168));
 sky130_fd_sc_hd__a41o_1 c293 (.A1(net1124),
    .A2(net48),
    .A3(net1104),
    .A4(net1118),
    .B1(net611),
    .X(net169));
 sky130_fd_sc_hd__mux4_1 c294 (.A0(net169),
    .A1(net165),
    .A2(net1086),
    .A3(net58),
    .S0(net132),
    .S1(clknet_1_0__leaf_net743),
    .X(net170));
 sky130_fd_sc_hd__mux4_1 c295 (.A0(net150),
    .A1(net1109),
    .A2(net161),
    .A3(net166),
    .S0(net1090),
    .S1(net1133),
    .X(net171));
 sky130_fd_sc_hd__a41o_2 c296 (.A1(net1071),
    .A2(net166),
    .A3(net883),
    .A4(net1111),
    .B1(net611),
    .X(net172));
 sky130_fd_sc_hd__mux4_1 c297 (.A0(net40),
    .A1(net169),
    .A2(net49),
    .A3(net883),
    .S0(net1028),
    .S1(net1054),
    .X(net173));
 sky130_fd_sc_hd__mux4_1 c298 (.A0(net895),
    .A1(clknet_1_0__leaf_net164),
    .A2(net172),
    .A3(net1090),
    .S0(net709),
    .S1(net752),
    .X(net174));
 sky130_fd_sc_hd__mux4_1 c299 (.A0(net153),
    .A1(net150),
    .A2(net172),
    .A3(net751),
    .S0(net752),
    .S1(net753),
    .X(net175));
 sky130_fd_sc_hd__mux4_1 c300 (.A0(clknet_1_1__leaf_net164),
    .A1(net172),
    .A2(net1112),
    .A3(net708),
    .S0(net748),
    .S1(net752),
    .X(net176));
 sky130_fd_sc_hd__mux4_1 c301 (.A0(net46),
    .A1(net48),
    .A2(net172),
    .A3(net1070),
    .S0(net974),
    .S1(net1080),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 c302 (.A0(clknet_1_0__leaf_net164),
    .A1(net172),
    .A2(net873),
    .A3(net1050),
    .S0(net1112),
    .S1(net753),
    .X(net178));
 sky130_fd_sc_hd__sdfbbn_1 c303 (.CLK_N(clknet_leaf_43_clk),
    .D(net49),
    .RESET_B(net172),
    .SCD(net161),
    .SCE(net691),
    .SET_B(net700),
    .Q(net180),
    .Q_N(net179));
 sky130_fd_sc_hd__mux4_2 c304 (.A0(net180),
    .A1(net52),
    .A2(net627),
    .A3(net629),
    .S0(clknet_1_0__leaf_net705),
    .S1(net749),
    .X(net181));
 sky130_fd_sc_hd__mux4_1 c305 (.A0(net172),
    .A1(net1122),
    .A2(net709),
    .A3(net1171),
    .S0(net754),
    .S1(net1140),
    .X(net182));
 sky130_fd_sc_hd__mux4_1 c306 (.A0(clknet_1_0__leaf_net181),
    .A1(net1053),
    .A2(net179),
    .A3(net605),
    .S0(net1128),
    .S1(net708),
    .X(net183));
 sky130_fd_sc_hd__mux4_1 c307 (.A0(net172),
    .A1(clknet_1_1__leaf_net183),
    .A2(net153),
    .A3(net605),
    .S0(net618),
    .S1(net754),
    .X(net184));
 sky130_fd_sc_hd__mux4_1 c308 (.A0(net925),
    .A1(net54),
    .A2(net1112),
    .A3(clknet_1_0__leaf_net704),
    .S0(clknet_1_0__leaf_net743),
    .S1(net750),
    .X(net185));
 sky130_fd_sc_hd__mux4_1 c309 (.A0(clknet_1_1__leaf_net164),
    .A1(net1093),
    .A2(net1110),
    .A3(net137),
    .S0(net1129),
    .S1(net1080),
    .X(net186));
 sky130_fd_sc_hd__sdfbbp_1 c310 (.CLK(clknet_leaf_43_clk),
    .D(net914),
    .RESET_B(net180),
    .SCD(net1055),
    .SCE(net1093),
    .SET_B(net1087),
    .Q(net188),
    .Q_N(net187));
 sky130_fd_sc_hd__a41o_1 c311 (.A1(net925),
    .A2(net914),
    .A3(clknet_1_0__leaf_net185),
    .A4(net750),
    .B1(net752),
    .X(net189));
 sky130_fd_sc_hd__mux4_1 c312 (.A0(net169),
    .A1(net907),
    .A2(net1107),
    .A3(net911),
    .S0(net1054),
    .S1(net914),
    .X(net190));
 sky130_fd_sc_hd__mux4_1 c313 (.A0(net898),
    .A1(net915),
    .A2(clknet_1_0__leaf_net704),
    .A3(clknet_1_0__leaf_net744),
    .S0(net751),
    .S1(net760),
    .X(net1002));
 sky130_fd_sc_hd__mux4_1 c314 (.A0(net136),
    .A1(net916),
    .A2(net1068),
    .A3(net986),
    .S0(net58),
    .S1(clknet_1_0__leaf_net185),
    .X(net191));
 sky130_fd_sc_hd__mux4_1 c315 (.A0(clknet_1_0__leaf_net191),
    .A1(net1073),
    .A2(net922),
    .A3(clknet_1_0__leaf_net183),
    .S0(net629),
    .S1(net759),
    .X(net192));
 sky130_fd_sc_hd__mux4_1 c316 (.A0(net897),
    .A1(net188),
    .A2(net907),
    .A3(clknet_1_0__leaf_net185),
    .S0(net165),
    .S1(clknet_1_0__leaf_net704),
    .X(net193));
 sky130_fd_sc_hd__sdfbbn_2 c317 (.CLK_N(clknet_leaf_44_clk),
    .D(clknet_1_1__leaf_net185),
    .RESET_B(clknet_1_0__leaf_net1002),
    .SCD(net1055),
    .SCE(net78),
    .SET_B(net757),
    .Q(net1009),
    .Q_N(net194));
 sky130_fd_sc_hd__mux4_2 c318 (.A0(net881),
    .A1(net1009),
    .A2(net612),
    .A3(net1080),
    .S0(net757),
    .S1(net759),
    .X(net195));
 sky130_fd_sc_hd__mux4_1 c319 (.A0(net898),
    .A1(net194),
    .A2(net37),
    .A3(net897),
    .S0(net1080),
    .S1(net1141),
    .X(net196));
 sky130_fd_sc_hd__mux4_1 c320 (.A0(net72),
    .A1(clknet_1_0__leaf_net189),
    .A2(net1009),
    .A3(net187),
    .S0(net141),
    .S1(net1064),
    .X(net197));
 sky130_fd_sc_hd__mux4_1 c321 (.A0(net907),
    .A1(net1055),
    .A2(clknet_1_0__leaf_net197),
    .A3(net1014),
    .S0(net760),
    .S1(net761),
    .X(net198));
 sky130_fd_sc_hd__mux4_1 c322 (.A0(net150),
    .A1(clknet_1_1__leaf_net185),
    .A2(net925),
    .A3(net1064),
    .S0(net1131),
    .S1(net762),
    .X(net199));
 sky130_fd_sc_hd__mux4_1 c323 (.A0(clknet_1_0__leaf_net183),
    .A1(clknet_1_0__leaf_net979),
    .A2(net890),
    .A3(clknet_1_1__leaf_net185),
    .S0(net1064),
    .S1(net757),
    .X(net200));
 sky130_fd_sc_hd__mux4_1 c324 (.A0(clknet_1_0__leaf_net197),
    .A1(net1064),
    .A2(clknet_1_0__leaf_net703),
    .A3(net760),
    .S0(net763),
    .S1(clknet_1_0__leaf_net764),
    .X(net201));
 sky130_fd_sc_hd__mux4_1 c325 (.A0(net152),
    .A1(net187),
    .A2(net1064),
    .A3(net194),
    .S0(net762),
    .S1(clknet_1_0__leaf_net765),
    .X(net996));
 sky130_fd_sc_hd__mux4_1 c326 (.A0(clknet_1_0__leaf_net996),
    .A1(net77),
    .A2(net1006),
    .A3(net194),
    .S0(net762),
    .S1(clknet_1_0__leaf_net764),
    .X(net202));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(net188),
    .A1(net150),
    .A2(clknet_1_0__leaf_net202),
    .A3(clknet_1_1__leaf_net191),
    .S0(net1126),
    .S1(clknet_1_0__leaf_net765),
    .X(net203));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(clknet_1_0__leaf_net202),
    .A1(net1107),
    .A2(clknet_1_0__leaf_net996),
    .A3(net1064),
    .S0(net1014),
    .S1(clknet_1_0__leaf_net703),
    .X(net204));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net1064),
    .A1(net165),
    .A2(clknet_1_0__leaf_net1002),
    .A3(clknet_1_0__leaf_net202),
    .S0(net691),
    .S1(clknet_1_0__leaf_net765),
    .X(net205));
 sky130_fd_sc_hd__mux4_1 c330 (.A0(clknet_1_1__leaf_net104),
    .A1(net1092),
    .A2(net916),
    .A3(net58),
    .S0(net1102),
    .S1(net890),
    .X(net206));
 sky130_fd_sc_hd__mux4_1 c331 (.A0(net941),
    .A1(net22),
    .A2(net172),
    .A3(net974),
    .S0(net719),
    .S1(clknet_1_0__leaf_net764),
    .X(net207));
 sky130_fd_sc_hd__mux4_1 c332 (.A0(net172),
    .A1(net1068),
    .A2(net871),
    .A3(net893),
    .S0(clknet_1_1__leaf_net635),
    .S1(clknet_1_1__leaf_net764),
    .X(net208));
 sky130_fd_sc_hd__mux4_1 c333 (.A0(clknet_1_1__leaf_net1002),
    .A1(net929),
    .A2(clknet_1_0__leaf_net206),
    .A3(net1014),
    .S0(net714),
    .S1(net763),
    .X(net209));
 sky130_fd_sc_hd__mux4_1 c334 (.A0(clknet_1_0__leaf_net206),
    .A1(clknet_1_0__leaf_net100),
    .A2(net1092),
    .A3(net163),
    .S0(net908),
    .S1(net761),
    .X(net210));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(clknet_1_1__leaf_net1002),
    .A1(net881),
    .A2(net605),
    .A3(net1014),
    .S0(clknet_1_1__leaf_net724),
    .S1(net731),
    .X(net211));
 sky130_fd_sc_hd__mux4_1 c336 (.A0(clknet_1_1__leaf_net88),
    .A1(net1064),
    .A2(clknet_1_1__leaf_net703),
    .A3(clknet_1_1__leaf_net726),
    .S0(net1077),
    .S1(clknet_1_1__leaf_net766),
    .X(net212));
 sky130_fd_sc_hd__mux4_2 c337 (.A0(net948),
    .A1(net77),
    .A2(net612),
    .A3(net631),
    .S0(net727),
    .S1(net1077),
    .X(net213));
 sky130_fd_sc_hd__mux4_1 c338 (.A0(net180),
    .A1(net1092),
    .A2(net213),
    .A3(clknet_1_0__leaf_net211),
    .S0(clknet_1_0__leaf_net996),
    .S1(net759),
    .X(net214));
 sky130_fd_sc_hd__mux4_1 c339 (.A0(net937),
    .A1(clknet_1_0__leaf_net211),
    .A2(net1006),
    .A3(net213),
    .S0(net920),
    .S1(net1131),
    .X(net215));
 sky130_fd_sc_hd__mux4_1 c340 (.A0(net141),
    .A1(net35),
    .A2(clknet_1_0__leaf_net215),
    .A3(net948),
    .S0(net597),
    .S1(clknet_1_0__leaf_net766),
    .X(net216));
 sky130_fd_sc_hd__mux4_1 c341 (.A0(net77),
    .A1(net1118),
    .A2(net671),
    .A3(clknet_1_0__leaf_net704),
    .S0(net713),
    .S1(net763),
    .X(net217));
 sky130_fd_sc_hd__mux4_1 c342 (.A0(net948),
    .A1(net938),
    .A2(net917),
    .A3(clknet_1_1__leaf_net100),
    .S0(net179),
    .S1(clknet_1_0__leaf_net766),
    .X(net990));
 sky130_fd_sc_hd__mux4_1 c343 (.A0(net1106),
    .A1(net1057),
    .A2(clknet_1_1__leaf_net88),
    .A3(clknet_1_0__leaf_net214),
    .S0(net605),
    .S1(net1014),
    .X(net218));
 sky130_fd_sc_hd__mux4_1 c344 (.A0(net213),
    .A1(clknet_1_0__leaf_net214),
    .A2(net909),
    .A3(net1072),
    .S0(net921),
    .S1(net597),
    .X(net219));
 sky130_fd_sc_hd__mux4_1 c345 (.A0(clknet_1_1__leaf_net206),
    .A1(net1096),
    .A2(net1132),
    .A3(net631),
    .S0(net676),
    .S1(net769),
    .X(net220));
 sky130_fd_sc_hd__mux4_1 c346 (.A0(net40),
    .A1(clknet_1_1__leaf_net202),
    .A2(clknet_1_0__leaf_net217),
    .A3(clknet_1_1__leaf_net211),
    .S0(net52),
    .S1(net771),
    .X(net221));
 sky130_fd_sc_hd__mux4_1 c347 (.A0(clknet_1_1__leaf_net211),
    .A1(net1064),
    .A2(clknet_1_1__leaf_net88),
    .A3(clknet_1_1__leaf_net765),
    .S0(net770),
    .S1(net1007),
    .X(net222));
 sky130_fd_sc_hd__mux4_1 c348 (.A0(net954),
    .A1(clknet_1_0__leaf_net990),
    .A2(clknet_1_0__leaf_net1022),
    .A3(net759),
    .S0(net771),
    .S1(net1007),
    .X(net223));
 sky130_fd_sc_hd__mux4_1 c349 (.A0(clknet_1_1__leaf_net103),
    .A1(clknet_1_0__leaf_net211),
    .A2(clknet_1_0__leaf_net193),
    .A3(clknet_1_0__leaf_net217),
    .S0(net676),
    .S1(net713),
    .X(net224));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(clknet_1_0__leaf_net217),
    .A1(net671),
    .A2(net676),
    .A3(net1001),
    .S0(net768),
    .S1(net770),
    .X(net225));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(clknet_1_1__leaf_net88),
    .A1(net213),
    .A2(clknet_1_0__leaf_net223),
    .A3(net631),
    .S0(clknet_1_0__leaf_net1022),
    .S1(net772),
    .X(net226));
 sky130_fd_sc_hd__mux4_1 c352 (.A0(clknet_1_1__leaf_net214),
    .A1(net962),
    .A2(net1072),
    .A3(net1102),
    .S0(net906),
    .S1(net763),
    .X(net227));
 sky130_fd_sc_hd__mux4_1 c353 (.A0(net143),
    .A1(net167),
    .A2(net78),
    .A3(net962),
    .S0(net691),
    .S1(net1077),
    .X(net228));
 sky130_fd_sc_hd__mux4_1 c354 (.A0(net228),
    .A1(net36),
    .A2(net940),
    .A3(clknet_1_1__leaf_net990),
    .S0(net736),
    .S1(clknet_1_1__leaf_net764),
    .X(net229));
 sky130_fd_sc_hd__mux4_1 c355 (.A0(net916),
    .A1(net3),
    .A2(clknet_1_1__leaf_net82),
    .A3(net166),
    .S0(net940),
    .S1(net735),
    .X(net230));
 sky130_fd_sc_hd__mux4_1 c356 (.A0(net228),
    .A1(net934),
    .A2(net966),
    .A3(net1023),
    .S0(net984),
    .S1(net676),
    .X(net231));
 sky130_fd_sc_hd__mux4_1 c357 (.A0(net0),
    .A1(clknet_1_1__leaf_net1002),
    .A2(net929),
    .A3(net741),
    .S0(net760),
    .S1(clknet_1_1__leaf_net764),
    .X(net232));
 sky130_fd_sc_hd__mux4_1 c358 (.A0(net1035),
    .A1(clknet_1_0__leaf_net232),
    .A2(net1110),
    .A3(net938),
    .S0(net997),
    .S1(net676),
    .X(net233));
 sky130_fd_sc_hd__mux4_1 c359 (.A0(net959),
    .A1(clknet_1_0__leaf_net233),
    .A2(net1023),
    .A3(clknet_1_0__leaf_net637),
    .S0(clknet_1_1__leaf_net705),
    .S1(net1077),
    .X(net234));
 sky130_fd_sc_hd__mux4_1 c360 (.A0(clknet_1_0__leaf_net232),
    .A1(net938),
    .A2(net3),
    .A3(net759),
    .S0(clknet_1_1__leaf_net766),
    .S1(net1013),
    .X(net235));
 sky130_fd_sc_hd__mux4_1 c361 (.A0(net929),
    .A1(net904),
    .A2(net1070),
    .A3(net961),
    .S0(net934),
    .S1(net721),
    .X(net1020));
 sky130_fd_sc_hd__mux4_1 c362 (.A0(net966),
    .A1(clknet_1_0__leaf_net113),
    .A2(net962),
    .A3(net633),
    .S0(net711),
    .S1(net995),
    .X(net236));
 sky130_fd_sc_hd__mux4_1 c363 (.A0(net938),
    .A1(clknet_1_1__leaf_net232),
    .A2(net1004),
    .A3(net672),
    .S0(net736),
    .S1(net1007),
    .X(net237));
 sky130_fd_sc_hd__mux4_1 c364 (.A0(net237),
    .A1(net1087),
    .A2(net734),
    .A3(net747),
    .S0(net763),
    .S1(net767),
    .X(net238));
 sky130_fd_sc_hd__mux4_1 c365 (.A0(clknet_1_0__leaf_net233),
    .A1(clknet_1_1__leaf_net214),
    .A2(net916),
    .A3(net881),
    .S0(net1033),
    .S1(net672),
    .X(net239));
 sky130_fd_sc_hd__mux4_1 c366 (.A0(clknet_1_1__leaf_net211),
    .A1(clknet_1_1__leaf_net113),
    .A2(net1126),
    .A3(net661),
    .S0(net760),
    .S1(net773),
    .X(net240));
 sky130_fd_sc_hd__mux4_1 c367 (.A0(net78),
    .A1(clknet_1_1__leaf_net217),
    .A2(net1033),
    .A3(net1036),
    .S0(net721),
    .S1(net1075),
    .X(net241));
 sky130_fd_sc_hd__mux4_1 c368 (.A0(net3),
    .A1(net1009),
    .A2(net966),
    .A3(net676),
    .S0(net734),
    .S1(clknet_1_1__leaf_net766),
    .X(net242));
 sky130_fd_sc_hd__mux4_1 c369 (.A0(net927),
    .A1(clknet_1_1__leaf_net113),
    .A2(clknet_1_0__leaf_net637),
    .A3(net1036),
    .S0(net1075),
    .S1(net775),
    .X(net243));
 sky130_fd_sc_hd__mux4_1 c370 (.A0(net167),
    .A1(net1036),
    .A2(net988),
    .A3(net722),
    .S0(net1075),
    .S1(net775),
    .X(net1029));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(clknet_1_1__leaf_net82),
    .A1(net1079),
    .A2(net720),
    .A3(net1077),
    .S0(net1075),
    .S1(net776),
    .X(net244));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net73),
    .A1(clknet_1_0__leaf_net241),
    .A2(clknet_1_1__leaf_net211),
    .A3(net228),
    .S0(net36),
    .S1(net775),
    .X(net245));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net244),
    .A1(clknet_1_1__leaf_net233),
    .A2(net1029),
    .A3(net661),
    .S0(net775),
    .S1(net777),
    .X(net246));
 sky130_fd_sc_hd__a41o_2 c396 (.A1(net144),
    .A2(net1123),
    .A3(net1091),
    .A4(net38),
    .B1(net1094),
    .X(net247));
 sky130_fd_sc_hd__sdfbbn_1 c397 (.CLK_N(clknet_leaf_7_clk),
    .D(net1056),
    .RESET_B(net1104),
    .SCD(net1108),
    .SCE(net1050),
    .SET_B(net1165),
    .Q(net249),
    .Q_N(net248));
 sky130_fd_sc_hd__a41o_1 c398 (.A1(net1049),
    .A2(net151),
    .A3(net149),
    .A4(net1124),
    .B1(net1082),
    .X(net250));
 sky130_fd_sc_hd__sdfbbp_1 c399 (.CLK(clknet_leaf_7_clk),
    .D(net1074),
    .RESET_B(net1094),
    .SCD(net1050),
    .SCE(net1082),
    .SET_B(clknet_1_1__leaf_net744),
    .Q(net252),
    .Q_N(net251));
 sky130_fd_sc_hd__sdfbbn_1 c400 (.CLK_N(clknet_leaf_7_clk),
    .D(net1049),
    .RESET_B(net1050),
    .SCD(net879),
    .SCE(net698),
    .SET_B(net1135),
    .Q(net254),
    .Q_N(net253));
 sky130_fd_sc_hd__a41o_1 c401 (.A1(net974),
    .A2(net1106),
    .A3(net610),
    .A4(clknet_1_0__leaf_net745),
    .B1(net746),
    .X(net255));
 sky130_fd_sc_hd__a41o_1 c402 (.A1(clknet_1_0__leaf_net255),
    .A2(net133),
    .A3(net1116),
    .A4(net616),
    .B1(net1082),
    .X(net256));
 sky130_fd_sc_hd__mux4_1 c403 (.A0(clknet_1_0__leaf_net256),
    .A1(net870),
    .A2(net248),
    .A3(net616),
    .S0(clknet_1_0__leaf_net745),
    .S1(net1134),
    .X(net257));
 sky130_fd_sc_hd__sdfbbn_1 c404 (.CLK_N(clknet_leaf_9_clk),
    .D(net252),
    .RESET_B(net1158),
    .SCD(net1094),
    .SCE(net135),
    .SET_B(net1049),
    .Q(net259),
    .Q_N(net258));
 sky130_fd_sc_hd__a41o_2 c405 (.A1(net254),
    .A2(net1123),
    .A3(net248),
    .A4(net1106),
    .B1(net1094),
    .X(net260));
 sky130_fd_sc_hd__a41o_1 c406 (.A1(clknet_1_0__leaf_net255),
    .A2(clknet_1_0__leaf_net256),
    .A3(net1092),
    .A4(net700),
    .B1(net1174),
    .X(net261));
 sky130_fd_sc_hd__sdfbbp_1 c407 (.CLK(clknet_leaf_8_clk),
    .D(net260),
    .RESET_B(net258),
    .SCD(net253),
    .SCE(clknet_1_0__leaf_net257),
    .SET_B(net1147),
    .Q(net263),
    .Q_N(net262));
 sky130_fd_sc_hd__sdfbbn_2 c408 (.CLK_N(clknet_leaf_9_clk),
    .D(clknet_1_1__leaf_net256),
    .RESET_B(clknet_1_1__leaf_net257),
    .SCD(net262),
    .SCE(net1051),
    .SET_B(net1115),
    .Q(net265),
    .Q_N(net264));
 sky130_fd_sc_hd__sdfbbn_2 c409 (.CLK_N(clknet_leaf_10_clk),
    .D(net1155),
    .RESET_B(net260),
    .SCD(net38),
    .SCE(net1049),
    .SET_B(clknet_1_0__leaf_net261),
    .Q(net267),
    .Q_N(net266));
 sky130_fd_sc_hd__mux4_2 c410 (.A0(net265),
    .A1(net1107),
    .A2(net142),
    .A3(net1069),
    .S0(net253),
    .S1(net616),
    .X(net268));
 sky130_fd_sc_hd__a41o_1 c411 (.A1(net263),
    .A2(net1074),
    .A3(net264),
    .A4(clknet_1_0__leaf_net256),
    .B1(net258),
    .X(net269));
 sky130_fd_sc_hd__mux4_1 c412 (.A0(net873),
    .A1(clknet_1_0__leaf_net255),
    .A2(net268),
    .A3(net260),
    .S0(net1050),
    .S1(clknet_1_0__leaf_net256),
    .X(net270));
 sky130_fd_sc_hd__mux4_1 c413 (.A0(net268),
    .A1(net144),
    .A2(net249),
    .A3(net262),
    .S0(clknet_1_0__leaf_net257),
    .S1(net1093),
    .X(net271));
 sky130_fd_sc_hd__mux4_1 c414 (.A0(net23),
    .A1(net268),
    .A2(net264),
    .A3(clknet_1_0__leaf_net269),
    .S0(net1136),
    .S1(net779),
    .X(net272));
 sky130_fd_sc_hd__sdfbbp_1 c415 (.CLK(clknet_leaf_7_clk),
    .D(net260),
    .RESET_B(net268),
    .SCD(clknet_1_0__leaf_net269),
    .SCE(net1163),
    .SET_B(net1143),
    .Q(net274),
    .Q_N(net273));
 sky130_fd_sc_hd__mux4_1 c416 (.A0(net1091),
    .A1(clknet_1_0__leaf_net261),
    .A2(net260),
    .A3(net266),
    .S0(net273),
    .S1(net781),
    .X(net275));
 sky130_fd_sc_hd__mux4_1 c417 (.A0(net268),
    .A1(net266),
    .A2(net1049),
    .A3(net273),
    .S0(net616),
    .S1(net780),
    .X(net276));
 sky130_fd_sc_hd__mux4_1 c418 (.A0(net870),
    .A1(net46),
    .A2(net1053),
    .A3(net1126),
    .S0(clknet_1_0__leaf_net703),
    .S1(net756),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 c419 (.A0(net879),
    .A1(net165),
    .A2(net1054),
    .A3(net46),
    .S0(net1116),
    .S1(clknet_1_0__leaf_net745),
    .X(net278));
 sky130_fd_sc_hd__mux4_2 c420 (.A0(net893),
    .A1(clknet_1_0__leaf_net255),
    .A2(net904),
    .A3(net1053),
    .S0(net616),
    .S1(clknet_1_1__leaf_net782),
    .X(net279));
 sky130_fd_sc_hd__mux4_1 c421 (.A0(net165),
    .A1(clknet_1_1__leaf_net269),
    .A2(clknet_1_0__leaf_net279),
    .A3(net1120),
    .S0(net610),
    .S1(net752),
    .X(net280));
 sky130_fd_sc_hd__sdfbbn_1 c422 (.CLK_N(clknet_leaf_5_clk),
    .D(clknet_1_0__leaf_net261),
    .RESET_B(net273),
    .SCD(net904),
    .SCE(net709),
    .SET_B(clknet_1_0__leaf_net782),
    .Q(net282),
    .Q_N(net281));
 sky130_fd_sc_hd__mux4_1 c423 (.A0(net1108),
    .A1(clknet_1_0__leaf_net279),
    .A2(net1052),
    .A3(net161),
    .S0(net906),
    .S1(net903),
    .X(net283));
 sky130_fd_sc_hd__sdfbbn_2 c424 (.CLK_N(clknet_leaf_7_clk),
    .D(net895),
    .RESET_B(clknet_1_0__leaf_net279),
    .SCD(net262),
    .SCE(net614),
    .SET_B(clknet_1_0__leaf_net782),
    .Q(net285),
    .Q_N(net284));
 sky130_fd_sc_hd__mux4_1 c425 (.A0(net132),
    .A1(net284),
    .A2(net957),
    .A3(net903),
    .S0(net614),
    .S1(net756),
    .X(net286));
 sky130_fd_sc_hd__mux4_1 c426 (.A0(net282),
    .A1(clknet_1_0__leaf_net255),
    .A2(net904),
    .A3(net616),
    .S0(net709),
    .S1(clknet_1_1__leaf_net782),
    .X(net287));
 sky130_fd_sc_hd__sdfbbp_1 c427 (.CLK(clknet_leaf_3_clk),
    .D(clknet_1_0__leaf_net277),
    .RESET_B(net1091),
    .SCD(net957),
    .SCE(net614),
    .SET_B(net1145),
    .Q(net289),
    .Q_N(net288));
 sky130_fd_sc_hd__a41o_1 c428 (.A1(net1110),
    .A2(net23),
    .A3(net288),
    .A4(net700),
    .B1(clknet_1_0__leaf_net782),
    .X(net290));
 sky130_fd_sc_hd__mux4_1 c429 (.A0(net898),
    .A1(net281),
    .A2(net251),
    .A3(clknet_1_0__leaf_net287),
    .S0(net1085),
    .S1(net605),
    .X(net291));
 sky130_fd_sc_hd__sdfbbn_1 c430 (.CLK_N(clknet_leaf_5_clk),
    .D(clknet_1_1__leaf_net269),
    .RESET_B(net1058),
    .SCD(net284),
    .SCE(clknet_1_0__leaf_net291),
    .SET_B(net1118),
    .Q(net293),
    .Q_N(net292));
 sky130_fd_sc_hd__mux4_1 c431 (.A0(net48),
    .A1(clknet_1_0__leaf_net277),
    .A2(net285),
    .A3(clknet_1_0__leaf_net279),
    .S0(net292),
    .S1(clknet_1_0__leaf_net783),
    .X(net294));
 sky130_fd_sc_hd__mux4_1 c432 (.A0(net47),
    .A1(net248),
    .A2(clknet_1_0__leaf_net290),
    .A3(net1163),
    .S0(clknet_1_0__leaf_net783),
    .S1(clknet_1_0__leaf_net784),
    .X(net295));
 sky130_fd_sc_hd__mux4_1 c433 (.A0(clknet_1_1__leaf_net287),
    .A1(net292),
    .A2(net288),
    .A3(net1071),
    .S0(net1116),
    .S1(net785),
    .X(net296));
 sky130_fd_sc_hd__mux4_1 c434 (.A0(net957),
    .A1(clknet_1_0__leaf_net296),
    .A2(clknet_1_0__leaf_net291),
    .A3(net49),
    .S0(clknet_1_0__leaf_net783),
    .S1(clknet_1_1__leaf_net784),
    .X(net297));
 sky130_fd_sc_hd__a41o_2 c435 (.A1(net1068),
    .A2(net292),
    .A3(net273),
    .A4(net605),
    .B1(net978),
    .X(net298));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(clknet_1_0__leaf_net290),
    .A1(clknet_1_0__leaf_net287),
    .A2(clknet_1_0__leaf_net979),
    .A3(net284),
    .S0(clknet_1_1__leaf_net784),
    .S1(net787),
    .X(net299));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(net298),
    .A1(net1127),
    .A2(net1055),
    .A3(clknet_1_0__leaf_net784),
    .S0(net787),
    .S1(net789),
    .X(net300));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(net293),
    .A1(net298),
    .A2(net284),
    .A3(clknet_1_0__leaf_net783),
    .S0(net786),
    .S1(net787),
    .X(net301));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net282),
    .A1(net298),
    .A2(clknet_1_0__leaf_net301),
    .S0(net756),
    .S1(net788),
    .X(net302));
 sky130_fd_sc_hd__mux4_2 c440 (.A0(net1110),
    .A1(net73),
    .A2(net298),
    .A3(net880),
    .S0(net691),
    .S1(net758),
    .X(net303));
 sky130_fd_sc_hd__mux4_1 c441 (.A0(net152),
    .A1(clknet_1_0__leaf_net1003),
    .A2(net35),
    .A3(net303),
    .S0(net752),
    .S1(net978),
    .X(net304));
 sky130_fd_sc_hd__mux4_1 c442 (.A0(net149),
    .A1(net188),
    .A2(net906),
    .A3(net974),
    .S0(net1093),
    .S1(net1137),
    .X(net305));
 sky130_fd_sc_hd__mux4_1 c443 (.A0(net267),
    .A1(net298),
    .A2(net264),
    .A3(net1065),
    .S0(net691),
    .S1(net790),
    .X(net306));
 sky130_fd_sc_hd__mux4_1 c444 (.A0(net1106),
    .A1(net911),
    .A2(net303),
    .A3(net1057),
    .S0(net790),
    .S1(net791),
    .X(net307));
 sky130_fd_sc_hd__mux4_1 c445 (.A0(net907),
    .A1(net915),
    .A2(net927),
    .A3(clknet_1_0__leaf_net202),
    .S0(net1054),
    .S1(net792),
    .X(net308));
 sky130_fd_sc_hd__mux4_1 c446 (.A0(clknet_1_0__leaf_net301),
    .A1(net1100),
    .A2(net35),
    .A3(net754),
    .S0(net791),
    .S1(net792),
    .X(net309));
 sky130_fd_sc_hd__mux4_1 c447 (.A0(net306),
    .A1(net303),
    .A2(net905),
    .A3(net758),
    .S0(clknet_1_0__leaf_net783),
    .S1(net792),
    .X(net310));
 sky130_fd_sc_hd__mux4_1 c448 (.A0(net281),
    .A1(clknet_1_1__leaf_net197),
    .A2(net652),
    .A3(net706),
    .S0(net758),
    .S1(net786),
    .X(net311));
 sky130_fd_sc_hd__mux4_1 c449 (.A0(net957),
    .A1(net1068),
    .A2(net909),
    .A3(net1053),
    .S0(net1076),
    .S1(net1011),
    .X(net312));
 sky130_fd_sc_hd__mux4_1 c450 (.A0(net77),
    .A1(net37),
    .A2(clknet_1_1__leaf_net255),
    .A3(net312),
    .S0(net1109),
    .S1(net1076),
    .X(net313));
 sky130_fd_sc_hd__mux4_1 c451 (.A0(net1052),
    .A1(net903),
    .A2(net696),
    .A3(net789),
    .S0(net790),
    .S1(net794),
    .X(net314));
 sky130_fd_sc_hd__mux4_2 c452 (.A0(net73),
    .A1(net1091),
    .A2(net707),
    .A3(net757),
    .S0(net791),
    .S1(net793),
    .X(net315));
 sky130_fd_sc_hd__mux4_1 c453 (.A0(net298),
    .A1(clknet_1_0__leaf_net197),
    .A2(net315),
    .A3(clknet_1_0__leaf_net277),
    .S0(net621),
    .S1(clknet_1_0__leaf_net743),
    .X(net316));
 sky130_fd_sc_hd__mux4_1 c454 (.A0(net162),
    .A1(net55),
    .A2(clknet_1_1__leaf_net261),
    .A3(net315),
    .S0(net652),
    .S1(net796),
    .X(net317));
 sky130_fd_sc_hd__mux4_1 c455 (.A0(clknet_1_1__leaf_net189),
    .A1(net306),
    .A2(net267),
    .A3(net315),
    .S0(net1011),
    .S1(net798),
    .X(net318));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(net312),
    .A1(net621),
    .A2(net790),
    .A3(net796),
    .S0(net798),
    .S1(net1015),
    .X(net319));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(clknet_1_1__leaf_net296),
    .A1(net622),
    .A2(net652),
    .A3(net798),
    .S0(net1015),
    .S1(clknet_1_0__leaf_net800),
    .X(net320));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(net909),
    .A1(net898),
    .A2(net1071),
    .A3(net303),
    .S0(net49),
    .S1(clknet_1_0__leaf_net800),
    .X(net321));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net274),
    .A1(clknet_1_1__leaf_net301),
    .A3(net715),
    .S0(net788),
    .S1(net791),
    .X(net322));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(clknet_1_1__leaf_net290),
    .A1(clknet_1_0__leaf_net999),
    .A2(clknet_1_1__leaf_net745),
    .A3(net758),
    .S0(net761),
    .S1(net799),
    .X(net323));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net1064),
    .A1(net655),
    .A2(clknet_1_0__leaf_net999),
    .A3(net758),
    .S0(net788),
    .S1(clknet_1_0__leaf_net801),
    .X(net324));
 sky130_fd_sc_hd__mux4_1 c462 (.A0(net909),
    .A1(net263),
    .A2(net1072),
    .A3(clknet_1_0__leaf_net1022),
    .S0(clknet_1_0__leaf_net704),
    .S1(net796),
    .X(net325));
 sky130_fd_sc_hd__mux4_2 c463 (.A0(net213),
    .A1(net940),
    .A2(net263),
    .A3(net1082),
    .S0(net769),
    .S1(net1011),
    .X(net326));
 sky130_fd_sc_hd__mux4_1 c464 (.A0(clknet_1_0__leaf_net325),
    .A1(net618),
    .A2(clknet_1_0__leaf_net1022),
    .A3(clknet_1_1__leaf_net726),
    .S0(net767),
    .S1(net1011),
    .X(net327));
 sky130_fd_sc_hd__mux4_1 c465 (.A0(clknet_1_1__leaf_net193),
    .A1(clknet_1_0__leaf_net324),
    .A2(net213),
    .A3(net40),
    .S0(net1097),
    .S1(net794),
    .X(net328));
 sky130_fd_sc_hd__mux4_1 c466 (.A0(net274),
    .A1(clknet_1_0__leaf_net328),
    .A2(net1061),
    .A3(net718),
    .S0(net1076),
    .S1(net795),
    .X(net329));
 sky130_fd_sc_hd__mux4_1 c467 (.A0(clknet_1_1__leaf_net325),
    .A1(net1102),
    .A2(net274),
    .A3(clknet_1_1__leaf_net635),
    .S0(net1077),
    .S1(net761),
    .X(net330));
 sky130_fd_sc_hd__mux4_1 c468 (.A0(net273),
    .A1(net285),
    .A2(net871),
    .A3(net631),
    .S0(net761),
    .S1(clknet_1_0__leaf_net802),
    .X(net331));
 sky130_fd_sc_hd__mux4_1 c469 (.A0(clknet_1_1__leaf_net255),
    .A1(net909),
    .A2(net691),
    .A3(net1076),
    .S0(clknet_1_1__leaf_net802),
    .S1(net803),
    .X(net332));
 sky130_fd_sc_hd__mux4_1 c470 (.A0(clknet_1_1__leaf_net331),
    .A1(clknet_1_1__leaf_net202),
    .A2(net1099),
    .A3(clknet_1_0__leaf_net332),
    .S0(net1007),
    .S1(net804),
    .X(net333));
 sky130_fd_sc_hd__mux4_1 c471 (.A0(net941),
    .A1(clknet_1_0__leaf_net223),
    .A2(net882),
    .A3(net1078),
    .S0(net754),
    .S1(clknet_1_0__leaf_net802),
    .X(net334));
 sky130_fd_sc_hd__mux4_1 c472 (.A0(net22),
    .A1(net940),
    .A2(clknet_1_1__leaf_net88),
    .A3(net251),
    .S0(clknet_1_1__leaf_net703),
    .S1(net731),
    .X(net335));
 sky130_fd_sc_hd__sdfbbn_1 c473 (.CLK_N(clknet_leaf_29_clk),
    .D(clknet_1_1__leaf_net202),
    .RESET_B(net1049),
    .SCD(net1102),
    .SCE(net1012),
    .SET_B(clknet_1_0__leaf_net801),
    .Q(net971),
    .Q_N(net336));
 sky130_fd_sc_hd__mux4_1 c474 (.A0(clknet_1_1__leaf_net279),
    .A1(net909),
    .A2(net672),
    .A3(net712),
    .S0(clknet_1_1__leaf_net802),
    .S1(net804),
    .X(net337));
 sky130_fd_sc_hd__mux4_1 c475 (.A0(net326),
    .A1(net920),
    .A2(net658),
    .A3(clknet_1_0__leaf_net1022),
    .S0(net710),
    .S1(net797),
    .X(net338));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(net940),
    .A1(net618),
    .A2(net631),
    .A3(net697),
    .S0(net768),
    .S1(clknet_1_0__leaf_net802),
    .X(net1000));
 sky130_fd_sc_hd__mux4_1 c477 (.A0(clknet_1_1__leaf_net332),
    .A1(net74),
    .A2(net326),
    .A3(net640),
    .S0(net799),
    .S1(net985),
    .X(net339));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(clknet_1_0__leaf_net331),
    .A1(clknet_1_0__leaf_net990),
    .A2(net1014),
    .A3(net663),
    .S0(net805),
    .S1(net807),
    .X(net340));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(net336),
    .A1(clknet_1_0__leaf_net1000),
    .A2(net663),
    .A3(net717),
    .S0(net721),
    .S1(net727),
    .X(net341));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(clknet_1_1__leaf_net223),
    .A1(net326),
    .A2(clknet_1_0__leaf_net341),
    .A3(net163),
    .S0(clknet_1_0__leaf_net328),
    .S1(net795),
    .X(net342));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net24),
    .A1(clknet_1_0__leaf_net225),
    .A2(clknet_1_0__leaf_net340),
    .A3(net137),
    .S0(net48),
    .S1(clknet_1_0__leaf_net341),
    .X(net343));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(clknet_1_1__leaf_net341),
    .A1(net1049),
    .A2(clknet_1_0__leaf_net340),
    .A3(net803),
    .S0(net806),
    .S1(net808),
    .X(net344));
 sky130_fd_sc_hd__a41o_1 c483 (.A1(net1102),
    .A2(net640),
    .A3(net663),
    .A4(net975),
    .B1(net808),
    .X(net345));
 sky130_fd_sc_hd__mux4_1 c484 (.A0(net1114),
    .A1(net962),
    .A2(net1008),
    .A3(net619),
    .S0(net722),
    .S1(clknet_1_1__leaf_net765),
    .X(net346));
 sky130_fd_sc_hd__mux4_1 c485 (.A0(clknet_1_1__leaf_net113),
    .A1(net959),
    .A2(net940),
    .A3(clknet_1_1__leaf_net279),
    .S0(net1004),
    .S1(net776),
    .X(net347));
 sky130_fd_sc_hd__mux4_1 c486 (.A0(clknet_1_1__leaf_net112),
    .A1(clknet_1_1__leaf_net217),
    .A2(net871),
    .A3(net682),
    .S0(net735),
    .S1(net778),
    .X(net348));
 sky130_fd_sc_hd__mux4_2 c487 (.A0(net904),
    .A1(net920),
    .A2(net1098),
    .A3(net1004),
    .S0(net719),
    .S1(net1075),
    .X(net349));
 sky130_fd_sc_hd__mux4_1 c488 (.A0(clknet_1_1__leaf_net346),
    .A1(clknet_1_1__leaf_net112),
    .A2(net641),
    .A3(net740),
    .S0(net774),
    .S1(net1015),
    .X(net350));
 sky130_fd_sc_hd__mux4_1 c489 (.A0(net902),
    .A1(clknet_1_1__leaf_net987),
    .A2(net662),
    .A3(net720),
    .S0(net741),
    .S1(net778),
    .X(net351));
 sky130_fd_sc_hd__mux4_2 c490 (.A0(net1102),
    .A1(net36),
    .A2(net735),
    .A3(net748),
    .S0(net763),
    .S1(net1005),
    .X(net352));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(net282),
    .A1(clknet_1_0__leaf_net346),
    .A2(net662),
    .A3(net664),
    .S0(net747),
    .S1(net808),
    .X(net353));
 sky130_fd_sc_hd__mux4_1 c492 (.A0(net960),
    .A1(net143),
    .A2(clknet_1_1__leaf_net261),
    .A3(net352),
    .S0(net641),
    .S1(net741),
    .X(net354));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(net289),
    .A1(clknet_1_1__leaf_net979),
    .A2(net900),
    .A3(net736),
    .S0(net748),
    .S1(net776),
    .X(net355));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(clknet_1_1__leaf_net112),
    .A1(net352),
    .A2(net345),
    .A3(clknet_1_1__leaf_net979),
    .S0(net1077),
    .S1(net754),
    .X(net356));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(net350),
    .A1(net353),
    .A2(net315),
    .A3(net959),
    .S0(net1081),
    .S1(net741),
    .X(net357));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(net1004),
    .A1(net754),
    .A2(net1005),
    .A3(net1075),
    .S0(clknet_1_1__leaf_net782),
    .S1(net809),
    .X(net358));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(clknet_1_1__leaf_net83),
    .A1(clknet_1_1__leaf_net979),
    .A2(net664),
    .A3(net733),
    .S0(net1075),
    .S1(net797),
    .X(net359));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(clknet_1_1__leaf_net279),
    .A1(net348),
    .A2(clknet_1_1__leaf_net340),
    .A3(net949),
    .S0(net773),
    .S1(net985),
    .X(net360));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(net358),
    .A1(net1021),
    .A2(net59),
    .A3(net922),
    .S0(net629),
    .S1(net810),
    .X(net361));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(net162),
    .A1(net940),
    .A2(net1058),
    .A3(clknet_1_1__leaf_net637),
    .S0(net776),
    .S1(net810),
    .X(net362));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(net940),
    .A1(clknet_1_1__leaf_net88),
    .A2(net959),
    .A3(net1004),
    .S0(net749),
    .S1(net810),
    .X(net363));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(net936),
    .A1(net1101),
    .A2(net882),
    .A3(net722),
    .S0(net736),
    .S1(net1010),
    .X(net364));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(net36),
    .A1(net960),
    .A2(net739),
    .A3(clknet_1_1__leaf_net801),
    .S0(net809),
    .S1(net1010),
    .X(net365));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(clknet_1_1__leaf_net217),
    .A1(net263),
    .A2(net138),
    .A3(net777),
    .S0(net809),
    .S1(net812),
    .X(net998));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(net289),
    .A1(net364),
    .A2(clknet_1_1__leaf_net987),
    .A3(net665),
    .S0(net711),
    .S1(net812),
    .X(net366));
 sky130_fd_sc_hd__sdfbbp_1 c528 (.CLK(clknet_leaf_9_clk),
    .D(net1057),
    .RESET_B(clknet_1_1__leaf_net257),
    .SCD(net39),
    .SCE(net1115),
    .SET_B(net779),
    .Q(net368),
    .Q_N(net367));
 sky130_fd_sc_hd__a41o_1 c529 (.A1(net145),
    .A2(net249),
    .A3(net1088),
    .A4(net1058),
    .B1(net1069),
    .X(net369));
 sky130_fd_sc_hd__sdfbbn_1 c530 (.CLK_N(clknet_leaf_9_clk),
    .D(net153),
    .RESET_B(net1069),
    .SCD(net1100),
    .SCE(net253),
    .SET_B(net1051),
    .Q(net371),
    .Q_N(net370));
 sky130_fd_sc_hd__mux4_1 c531 (.A0(net259),
    .A1(net267),
    .A2(net1097),
    .A3(clknet_1_0__leaf_net261),
    .S0(net1115),
    .S1(net780),
    .X(net372));
 sky130_fd_sc_hd__a41o_2 c532 (.A1(net136),
    .A2(net254),
    .A3(net1073),
    .A4(net699),
    .B1(net1080),
    .X(net373));
 sky130_fd_sc_hd__sdfbbn_1 c533 (.CLK_N(clknet_leaf_9_clk),
    .D(net1127),
    .RESET_B(net1051),
    .SCD(net28),
    .SCE(net600),
    .SET_B(net1082),
    .Q(net991),
    .Q_N(net374));
 sky130_fd_sc_hd__sdfbbp_1 c534 (.CLK(clknet_leaf_11_clk),
    .D(net268),
    .RESET_B(net974),
    .SCD(net373),
    .SCE(clknet_1_1__leaf_net256),
    .SET_B(net1146),
    .Q(net376),
    .Q_N(net375));
 sky130_fd_sc_hd__a41o_4 c535 (.A1(net260),
    .A2(net1104),
    .A3(net1115),
    .A4(net779),
    .B1(net814),
    .X(net377));
 sky130_fd_sc_hd__mux4_1 c536 (.A0(net374),
    .A1(net377),
    .A2(net373),
    .A3(net1056),
    .S0(net1115),
    .S1(net616),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 c537 (.A0(net876),
    .A1(net377),
    .A2(net1056),
    .A3(net1115),
    .S0(net600),
    .S1(net780),
    .X(net379));
 sky130_fd_sc_hd__a41o_1 c538 (.A1(net377),
    .A2(net1100),
    .A3(net367),
    .A4(net600),
    .B1(net781),
    .X(net380));
 sky130_fd_sc_hd__sdfbbn_1 c539 (.CLK_N(clknet_leaf_10_clk),
    .D(net377),
    .RESET_B(net1069),
    .SCD(net39),
    .SCE(net1108),
    .SET_B(net380),
    .Q(net382),
    .Q_N(net381));
 sky130_fd_sc_hd__mux4_1 c540 (.A0(net368),
    .A1(net373),
    .A2(net1105),
    .A3(net1106),
    .S0(net28),
    .S1(net779),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 c541 (.A0(net145),
    .A1(net1123),
    .A2(net375),
    .A3(clknet_1_0__leaf_net999),
    .S0(net699),
    .S1(net815),
    .X(net384));
 sky130_fd_sc_hd__a41o_1 c542 (.A1(net1121),
    .A2(net1088),
    .A3(net259),
    .A4(net781),
    .B1(net816),
    .X(net385));
 sky130_fd_sc_hd__mux4_1 c543 (.A0(net380),
    .A1(net368),
    .A2(net1057),
    .A3(net1060),
    .S0(net385),
    .S1(net779),
    .X(net386));
 sky130_fd_sc_hd__a41o_1 c544 (.A1(net376),
    .A2(net381),
    .A3(net618),
    .A4(net816),
    .B1(clknet_1_0__leaf_net818),
    .X(net387));
 sky130_fd_sc_hd__mux4_1 c545 (.A0(net254),
    .A1(net1100),
    .A2(net373),
    .A3(net258),
    .S0(clknet_1_0__leaf_net387),
    .S1(clknet_1_0__leaf_net818),
    .X(net388));
 sky130_fd_sc_hd__a41o_1 c546 (.A1(net148),
    .A2(net385),
    .A3(clknet_1_1__leaf_net387),
    .A4(net817),
    .B1(clknet_1_0__leaf_net818),
    .X(net389));
 sky130_fd_sc_hd__a41o_1 c547 (.A1(net29),
    .A2(net1127),
    .A3(net381),
    .A4(clknet_1_1__leaf_net389),
    .B1(clknet_1_0__leaf_net818),
    .X(net390));
 sky130_fd_sc_hd__mux4_1 c548 (.A0(clknet_1_1__leaf_net256),
    .A1(clknet_1_1__leaf_net389),
    .A2(net382),
    .A3(net1117),
    .S0(clknet_1_0__leaf_net818),
    .S1(clknet_1_0__leaf_net819),
    .X(net391));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(clknet_1_1__leaf_net257),
    .A1(clknet_1_0__leaf_net387),
    .A2(clknet_1_0__leaf_net389),
    .A3(net370),
    .S0(net373),
    .S1(net142),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c550 (.A0(net376),
    .A1(net1121),
    .A2(net266),
    .A3(net284),
    .S0(net1120),
    .S1(net756),
    .X(net972));
 sky130_fd_sc_hd__mux4_1 c551 (.A0(net1062),
    .A1(net249),
    .A2(net284),
    .A3(net1128),
    .S0(net1137),
    .S1(clknet_1_0__leaf_net818),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 c552 (.A0(net162),
    .A1(net1073),
    .A2(net251),
    .A3(net1080),
    .S0(net756),
    .S1(clknet_1_0__leaf_net818),
    .X(net394));
 sky130_fd_sc_hd__mux4_1 c553 (.A0(clknet_1_0__leaf_net394),
    .A1(net49),
    .A2(net153),
    .A3(net1115),
    .S0(net700),
    .S1(clknet_1_0__leaf_net819),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 c554 (.A0(net252),
    .A1(net274),
    .A2(net1062),
    .A3(net1085),
    .S0(net752),
    .S1(clknet_1_0__leaf_net783),
    .X(net396));
 sky130_fd_sc_hd__mux4_2 c555 (.A0(net385),
    .A1(net163),
    .A2(net285),
    .A3(net267),
    .S0(net263),
    .S1(net1062),
    .X(net397));
 sky130_fd_sc_hd__mux4_2 c556 (.A0(clknet_1_0__leaf_net181),
    .A1(net385),
    .A2(net161),
    .A3(net614),
    .S0(clknet_1_1__leaf_net744),
    .S1(net816),
    .X(net398));
 sky130_fd_sc_hd__mux4_2 c557 (.A0(net895),
    .A1(net138),
    .A2(net1062),
    .A3(net903),
    .S0(net375),
    .S1(net1085),
    .X(net399));
 sky130_fd_sc_hd__mux4_1 c558 (.A0(net399),
    .A1(net65),
    .A2(net895),
    .A3(net135),
    .S0(net1123),
    .S1(clknet_1_0__leaf_net398),
    .X(net400));
 sky130_fd_sc_hd__mux4_1 c559 (.A0(net399),
    .A1(net376),
    .A2(clknet_1_0__leaf_net979),
    .A3(clknet_1_0__leaf_net396),
    .S0(net600),
    .S1(net1130),
    .X(net401));
 sky130_fd_sc_hd__mux4_1 c560 (.A0(net382),
    .A1(net1062),
    .A2(clknet_1_1__leaf_net394),
    .A3(net1106),
    .S0(net816),
    .S1(net821),
    .X(net402));
 sky130_fd_sc_hd__mux4_1 c561 (.A0(net1055),
    .A1(net1123),
    .A2(net266),
    .A3(net752),
    .S0(net817),
    .S1(net822),
    .X(net403));
 sky130_fd_sc_hd__a41o_1 c562 (.A1(net367),
    .A2(clknet_1_1__leaf_net181),
    .A3(net695),
    .A4(net813),
    .B1(net824),
    .X(net404));
 sky130_fd_sc_hd__mux4_1 c563 (.A0(clknet_1_1__leaf_net387),
    .A1(clknet_1_0__leaf_net400),
    .A2(net1062),
    .A3(clknet_1_1__leaf_net745),
    .S0(net822),
    .S1(net823),
    .X(net405));
 sky130_fd_sc_hd__mux4_2 c564 (.A0(clknet_1_1__leaf_net398),
    .A1(clknet_1_1__leaf_net181),
    .A2(net399),
    .A3(clknet_1_0__leaf_net820),
    .S0(net824),
    .S1(net825),
    .X(net406));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net1057),
    .A1(net1062),
    .A2(clknet_1_0__leaf_net406),
    .A3(clknet_1_0__leaf_net819),
    .S0(net823),
    .S1(net826),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(clknet_1_0__leaf_net406),
    .A1(clknet_1_0__leaf_net390),
    .A2(clknet_1_1__leaf_net404),
    .A3(clknet_1_1__leaf_net743),
    .S0(net787),
    .S1(net825),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c567 (.A0(clknet_1_1__leaf_net406),
    .A1(clknet_1_0__leaf_net651),
    .A2(net700),
    .A3(net785),
    .S0(net787),
    .S1(net821),
    .X(net409));
 sky130_fd_sc_hd__mux4_2 c568 (.A0(net249),
    .A1(net293),
    .A2(net1062),
    .A3(net817),
    .S0(net821),
    .S1(net827),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(clknet_1_1__leaf_net400),
    .A1(net136),
    .A2(clknet_1_0__leaf_net398),
    .A3(net410),
    .S0(net753),
    .S1(net817),
    .X(net411));
 sky130_fd_sc_hd__mux4_2 c570 (.A0(net410),
    .A1(clknet_1_1__leaf_net406),
    .A3(net822),
    .S0(net828),
    .S1(net829),
    .X(net651));
 sky130_fd_sc_hd__mux4_2 c571 (.A0(clknet_1_0__leaf_net398),
    .A1(clknet_1_0__leaf_net651),
    .A2(net978),
    .A3(net817),
    .S0(clknet_1_1__leaf_net819),
    .S1(net829),
    .X(net413));
 sky130_fd_sc_hd__mux4_1 c572 (.A0(clknet_1_0__leaf_net404),
    .A1(net991),
    .A2(net1057),
    .A3(net911),
    .S0(net752),
    .S1(net755),
    .X(net414));
 sky130_fd_sc_hd__mux4_1 c573 (.A0(clknet_1_1__leaf_net197),
    .A1(net1052),
    .A2(net927),
    .A3(net1097),
    .S0(clknet_1_1__leaf_net745),
    .S1(net752),
    .X(net415));
 sky130_fd_sc_hd__mux4_2 c574 (.A0(net399),
    .A1(net1102),
    .A2(net1078),
    .A3(net792),
    .S0(net815),
    .S1(net816),
    .X(net416));
 sky130_fd_sc_hd__mux4_1 c575 (.A0(net911),
    .A1(net303),
    .A2(net410),
    .A3(net1072),
    .S0(net656),
    .S1(net793),
    .X(net417));
 sky130_fd_sc_hd__mux4_1 c576 (.A0(net891),
    .A1(net315),
    .A2(net906),
    .A3(net1065),
    .S0(net656),
    .S1(net1159),
    .X(net418));
 sky130_fd_sc_hd__mux4_1 c577 (.A0(net922),
    .A1(net695),
    .A2(clknet_1_1__leaf_net800),
    .A3(net815),
    .S0(clknet_1_1__leaf_net820),
    .S1(net830),
    .X(net992));
 sky130_fd_sc_hd__mux4_1 c578 (.A0(net410),
    .A1(net1055),
    .A2(net1070),
    .A3(net927),
    .S0(net1173),
    .S1(clknet_1_1__leaf_net745),
    .X(net419));
 sky130_fd_sc_hd__mux4_1 c579 (.A0(net293),
    .A1(net1108),
    .A2(net1056),
    .A3(net262),
    .S0(net634),
    .S1(net815),
    .X(net420));
 sky130_fd_sc_hd__mux4_1 c580 (.A0(clknet_1_0__leaf_net296),
    .A1(net1099),
    .A2(clknet_1_1__leaf_net197),
    .A3(clknet_1_1__leaf_net819),
    .S0(net822),
    .S1(net828),
    .X(net421));
 sky130_fd_sc_hd__mux4_1 c581 (.A0(net267),
    .A1(net1053),
    .A2(net1097),
    .A3(net622),
    .S0(net829),
    .S1(net836),
    .X(net422));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(net422),
    .A1(net29),
    .A2(clknet_1_1__leaf_net197),
    .A3(net816),
    .S0(net832),
    .S1(net836),
    .X(net423));
 sky130_fd_sc_hd__mux4_1 c583 (.A0(net1108),
    .A1(net78),
    .A2(net600),
    .A3(net793),
    .S0(net1084),
    .S1(net837),
    .X(net424));
 sky130_fd_sc_hd__mux4_1 c584 (.A0(net29),
    .A1(net267),
    .A2(clknet_1_1__leaf_net800),
    .A3(net816),
    .S0(net827),
    .S1(net830),
    .X(net425));
 sky130_fd_sc_hd__mux4_1 c585 (.A0(clknet_1_1__leaf_net396),
    .A1(net900),
    .A2(net927),
    .A3(net187),
    .S0(net986),
    .S1(net1103),
    .X(net969));
 sky130_fd_sc_hd__mux4_1 c586 (.A0(net424),
    .A1(net416),
    .A2(net262),
    .A3(net251),
    .S0(clknet_1_1__leaf_net819),
    .S1(net837),
    .X(net426));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(clknet_1_0__leaf_net425),
    .A1(clknet_1_1__leaf_net296),
    .A2(net163),
    .A3(net1080),
    .S0(clknet_1_1__leaf_net783),
    .S1(net833),
    .X(net427));
 sky130_fd_sc_hd__mux4_1 c588 (.A0(net377),
    .A1(net424),
    .A2(net274),
    .A3(clknet_1_0__leaf_net393),
    .S0(net58),
    .S1(net817),
    .X(net428));
 sky130_fd_sc_hd__mux4_1 c589 (.A0(net49),
    .A1(clknet_1_1__leaf_net651),
    .A2(net982),
    .A3(net796),
    .S0(net836),
    .S1(net989),
    .X(net429));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(net974),
    .A1(clknet_1_1__leaf_net744),
    .A2(net816),
    .A3(net835),
    .S0(net837),
    .S1(net989),
    .X(net430));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(net399),
    .A1(net634),
    .A2(clknet_1_0__leaf_net801),
    .A3(net828),
    .S0(net1084),
    .S1(net837),
    .X(net431));
 sky130_fd_sc_hd__sdfbbn_1 c592 (.CLK_N(clknet_leaf_18_clk),
    .D(clknet_1_0__leaf_net431),
    .RESET_B(net1168),
    .SCD(net422),
    .SCE(net634),
    .SET_B(net793),
    .Q(net433),
    .Q_N(net432));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(clknet_1_1__leaf_net431),
    .A1(net432),
    .A2(net900),
    .A3(net989),
    .S0(clknet_1_0__leaf_net838),
    .S1(clknet_1_0__leaf_net839),
    .X(net434));
 sky130_fd_sc_hd__mux4_1 c594 (.A0(net374),
    .A1(clknet_1_0__leaf_net996),
    .A2(net1088),
    .A3(net695),
    .S0(net714),
    .S1(net834),
    .X(net435));
 sky130_fd_sc_hd__mux4_1 c595 (.A0(net274),
    .A1(clknet_1_1__leaf_net425),
    .A2(net949),
    .A3(net1089),
    .S0(net712),
    .S1(net806),
    .X(net436));
 sky130_fd_sc_hd__mux4_1 c596 (.A0(net298),
    .A1(net1056),
    .A2(clknet_1_0__leaf_net328),
    .A3(net1078),
    .S0(net790),
    .S1(net803),
    .X(net437));
 sky130_fd_sc_hd__mux4_1 c597 (.A0(net416),
    .A1(clknet_1_1__leaf_net202),
    .A2(clknet_1_0__leaf_net225),
    .A3(clknet_1_0__leaf_net990),
    .S0(net917),
    .S1(clknet_1_1__leaf_net703),
    .X(net438));
 sky130_fd_sc_hd__mux4_1 c598 (.A0(net436),
    .A1(net377),
    .A2(clknet_1_0__leaf_net990),
    .A3(net1118),
    .S0(net922),
    .S1(net826),
    .X(net439));
 sky130_fd_sc_hd__mux4_1 c599 (.A0(net397),
    .A1(clknet_1_0__leaf_net439),
    .A2(net880),
    .A3(net1049),
    .S0(clknet_1_1__leaf_net261),
    .S1(net804),
    .X(net440));
 sky130_fd_sc_hd__mux4_1 c600 (.A0(net48),
    .A1(clknet_1_0__leaf_net990),
    .A2(clknet_1_0__leaf_net340),
    .A3(net949),
    .S0(net285),
    .S1(clknet_1_0__leaf_net840),
    .X(net441));
 sky130_fd_sc_hd__mux4_1 c601 (.A0(clknet_1_0__leaf_net425),
    .A1(net974),
    .A2(net1103),
    .A3(net163),
    .S0(net941),
    .S1(net807),
    .X(net442));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(net1049),
    .A1(net433),
    .A2(clknet_1_0__leaf_net990),
    .A3(net941),
    .S0(net677),
    .S1(clknet_1_1__leaf_net818),
    .X(net443));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(clknet_1_1__leaf_net439),
    .A1(clknet_1_0__leaf_net992),
    .A2(net48),
    .A3(net714),
    .S0(net718),
    .S1(clknet_1_1__leaf_net801),
    .X(net444));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(clknet_1_1__leaf_net225),
    .A1(net345),
    .A2(clknet_1_0__leaf_net992),
    .A3(net949),
    .S0(net1099),
    .S1(net677),
    .X(net445));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(clknet_1_1__leaf_net290),
    .A1(net285),
    .A2(net1049),
    .A3(net677),
    .S0(net717),
    .S1(net831),
    .X(net446));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net163),
    .A1(net76),
    .A2(net41),
    .A3(net137),
    .S0(net1105),
    .S1(net1012),
    .X(net447));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(net1059),
    .A1(net658),
    .A2(net1040),
    .A3(net807),
    .S0(clknet_1_1__leaf_net818),
    .S1(clknet_1_1__leaf_net839),
    .X(net448));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net377),
    .A1(clknet_1_0__leaf_net435),
    .A2(net618),
    .A3(net788),
    .S0(net826),
    .S1(net842),
    .X(net449));
 sky130_fd_sc_hd__mux4_1 c609 (.A0(net416),
    .A1(net900),
    .A2(net660),
    .A3(net677),
    .S0(clknet_1_0__leaf_net840),
    .S1(net843),
    .X(net450));
 sky130_fd_sc_hd__mux4_2 c610 (.A0(net413),
    .A1(net73),
    .A2(clknet_1_0__leaf_net439),
    .A3(net1082),
    .S0(net772),
    .S1(net994),
    .X(net451));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net303),
    .A1(net949),
    .A2(net993),
    .A3(net978),
    .S0(clknet_1_1__leaf_net840),
    .S1(net843),
    .X(net452));
 sky130_fd_sc_hd__a41o_1 c612 (.A1(net906),
    .A2(net247),
    .A3(net660),
    .A4(net678),
    .B1(net1153),
    .X(net453));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(net41),
    .A1(clknet_1_1__leaf_net439),
    .A2(net1118),
    .A3(net678),
    .S0(net680),
    .S1(net841),
    .X(net454));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(net442),
    .A1(net162),
    .A2(net980),
    .A3(clknet_1_1__leaf_net802),
    .S0(clknet_1_1__leaf_net818),
    .S1(net843),
    .X(net455));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(clknet_1_1__leaf_net100),
    .A1(net882),
    .A2(net660),
    .A3(net680),
    .S0(net688),
    .S1(clknet_1_0__leaf_net840),
    .X(net456));
 sky130_fd_sc_hd__mux4_2 c616 (.A0(net263),
    .A1(net1021),
    .A2(net1106),
    .A3(net949),
    .S0(net1040),
    .S1(net1075),
    .X(net981));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(net1057),
    .A1(net1063),
    .A2(net917),
    .A3(net904),
    .S0(net981),
    .S1(clknet_1_1__leaf_net783),
    .X(net457));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(clknet_1_0__leaf_net365),
    .A1(net73),
    .A2(net162),
    .A3(net961),
    .S0(net927),
    .S1(net1078),
    .X(net458));
 sky130_fd_sc_hd__mux4_1 c619 (.A0(net349),
    .A1(net1072),
    .A2(clknet_1_0__leaf_net458),
    .A3(net682),
    .S0(clknet_1_1__leaf_net703),
    .S1(net827),
    .X(net459));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net900),
    .A1(net920),
    .A2(net1119),
    .A3(clknet_1_1__leaf_net361),
    .S0(clknet_1_1__leaf_net996),
    .S1(net1076),
    .X(net976));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(net1089),
    .A1(clknet_1_0__leaf_net365),
    .A2(clknet_1_1__leaf_net637),
    .A3(net661),
    .S0(net682),
    .S1(net994),
    .X(net460));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(clknet_1_0__leaf_net340),
    .A1(net352),
    .A2(net922),
    .A3(net1110),
    .S0(net1079),
    .S1(net1078),
    .X(net461));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(clknet_1_0__leaf_net361),
    .A1(clknet_1_1__leaf_net996),
    .A2(clknet_1_1__leaf_net990),
    .A3(net661),
    .S0(net694),
    .S1(clknet_1_1__leaf_net839),
    .X(net462));
 sky130_fd_sc_hd__mux4_1 c624 (.A0(net138),
    .A1(net927),
    .A2(clknet_1_0__leaf_net460),
    .A3(clknet_1_1__leaf_net291),
    .S0(clknet_1_1__leaf_net990),
    .S1(net749),
    .X(net463));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net917),
    .A1(net981),
    .A2(clknet_1_0__leaf_net460),
    .A3(net721),
    .S0(clknet_1_1__leaf_net839),
    .S1(net844),
    .X(net464));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net1109),
    .A1(net1101),
    .A2(net1097),
    .A3(net1081),
    .S0(net772),
    .S1(net799),
    .X(net465));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(net345),
    .A1(clknet_1_0__leaf_net464),
    .A2(clknet_1_0__leaf_net969),
    .A3(net432),
    .S0(net679),
    .S1(net749),
    .X(net466));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net1119),
    .A1(clknet_1_0__leaf_net976),
    .A2(net665),
    .A3(net694),
    .S0(net835),
    .S1(net989),
    .X(net467));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(net1072),
    .A1(net1089),
    .A2(net349),
    .A3(net1078),
    .S0(net1075),
    .S1(net799),
    .X(net468));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net468),
    .A1(net949),
    .A2(net465),
    .A3(clknet_1_0__leaf_net462),
    .S0(clknet_1_0__leaf_net458),
    .S1(net993),
    .X(net469));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net364),
    .A1(net882),
    .A2(net1109),
    .A3(net978),
    .S0(net797),
    .S1(net846),
    .X(net470));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(clknet_1_0__leaf_net462),
    .A1(net736),
    .A2(net1076),
    .A3(net773),
    .S0(net1075),
    .S1(net846),
    .X(net471));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(net465),
    .A1(net352),
    .A2(clknet_1_1__leaf_net462),
    .A3(net993),
    .S0(net772),
    .S1(net846),
    .X(net472));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net433),
    .A1(net1039),
    .A2(net986),
    .A3(net465),
    .S0(net1076),
    .S1(net845),
    .X(net473));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net473),
    .A1(net349),
    .A2(clknet_1_0__leaf_net361),
    .A3(net1101),
    .S0(clknet_1_1__leaf_net783),
    .S1(net975),
    .X(net474));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net906),
    .A1(net474),
    .A2(net473),
    .A3(clknet_1_1__leaf_net365),
    .S0(net694),
    .S1(net747),
    .X(net475));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net470),
    .A1(clknet_1_0__leaf_net970),
    .A2(net689),
    .A3(net721),
    .S0(net773),
    .S1(net827),
    .X(net476));
 sky130_fd_sc_hd__sdfbbp_1 c660 (.CLK(clknet_leaf_11_clk),
    .D(net1123),
    .RESET_B(net375),
    .SCD(net1073),
    .SCE(net1051),
    .SET_B(clknet_1_1__leaf_net999),
    .Q(net478),
    .Q_N(net477));
 sky130_fd_sc_hd__mux4_1 c661 (.A0(clknet_1_0__leaf_net389),
    .A1(net1051),
    .A2(net1127),
    .A3(net377),
    .S0(net1086),
    .S1(net1117),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c662 (.A0(net260),
    .A1(net1123),
    .A2(net477),
    .A3(net147),
    .S0(net38),
    .S1(net1082),
    .X(net480));
 sky130_fd_sc_hd__sdfbbn_1 c663 (.CLK_N(clknet_leaf_11_clk),
    .D(net368),
    .RESET_B(net1097),
    .SCD(clknet_1_0__leaf_net261),
    .SCE(net600),
    .SET_B(clknet_1_1__leaf_net999),
    .Q(net482),
    .Q_N(net481));
 sky130_fd_sc_hd__a41o_1 c664 (.A1(net1097),
    .A2(net481),
    .A3(net1051),
    .B1(clknet_1_0__leaf_net820),
    .X(net483));
 sky130_fd_sc_hd__sdfbbn_1 c665 (.CLK_N(clknet_leaf_11_clk),
    .D(net1160),
    .RESET_B(net1060),
    .SCD(net1053),
    .SCE(net260),
    .SET_B(net747),
    .Q(net485),
    .Q_N(net484));
 sky130_fd_sc_hd__sdfbbp_1 c666 (.CLK(clknet_leaf_11_clk),
    .D(net480),
    .RESET_B(net485),
    .SCD(net1051),
    .SCE(net1058),
    .SET_B(net1162),
    .Q(net487),
    .Q_N(net486));
 sky130_fd_sc_hd__a41o_1 c667 (.A1(net148),
    .A2(net1121),
    .A3(net486),
    .A4(net780),
    .B1(clknet_1_0__leaf_net818),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c668 (.A0(net1051),
    .A1(net480),
    .A2(net1097),
    .A3(net484),
    .S0(clknet_1_0__leaf_net488),
    .S1(net1083),
    .X(net489));
 sky130_fd_sc_hd__sdfbbn_1 c669 (.CLK_N(clknet_leaf_10_clk),
    .D(clknet_1_0__leaf_net261),
    .RESET_B(net367),
    .SCD(net370),
    .SCE(net781),
    .SET_B(net1154),
    .Q(net491),
    .Q_N(net490));
 sky130_fd_sc_hd__mux4_1 c670 (.A0(net487),
    .A1(net1106),
    .A2(clknet_1_0__leaf_net488),
    .A3(net147),
    .S0(net1051),
    .S1(net1083),
    .X(net492));
 sky130_fd_sc_hd__mux4_1 c671 (.A0(net268),
    .A1(net1117),
    .A2(net1115),
    .A3(net490),
    .S0(net609),
    .S1(clknet_1_1__leaf_net999),
    .X(net493));
 sky130_fd_sc_hd__sdfbbn_1 c672 (.CLK_N(clknet_leaf_12_clk),
    .D(clknet_1_0__leaf_net493),
    .RESET_B(net1157),
    .SCD(net1117),
    .SCE(net847),
    .SET_B(net1150),
    .Q(net495),
    .Q_N(net494));
 sky130_fd_sc_hd__sdfbbp_1 c673 (.CLK(clknet_leaf_11_clk),
    .D(net373),
    .RESET_B(net495),
    .SCD(net482),
    .SCE(net847),
    .SET_B(net848),
    .Q(net497),
    .Q_N(net496));
 sky130_fd_sc_hd__sdfbbn_1 c674 (.CLK_N(clknet_leaf_12_clk),
    .D(net497),
    .RESET_B(net1156),
    .SCD(net1058),
    .SCE(net1051),
    .SET_B(net1103),
    .Q(net499),
    .Q_N(net498));
 sky130_fd_sc_hd__mux4_2 c675 (.A0(net485),
    .A1(net495),
    .A2(net487),
    .A3(net499),
    .S0(net1121),
    .S1(net1083),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c676 (.A0(net380),
    .A1(net497),
    .A2(net477),
    .A3(net1108),
    .S0(clknet_1_0__leaf_net818),
    .S1(net1150),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c677 (.A0(clknet_1_1__leaf_net493),
    .A1(net499),
    .A2(net494),
    .A3(net1069),
    .S0(net847),
    .S1(net849),
    .X(net502));
 sky130_fd_sc_hd__a41o_1 c678 (.A1(net478),
    .A2(net498),
    .A3(clknet_1_1__leaf_net743),
    .A4(net847),
    .B1(net850),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c679 (.A0(net1087),
    .A1(clknet_1_0__leaf_net503),
    .A2(net498),
    .A3(net486),
    .S0(net608),
    .S1(net850),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c680 (.A0(clknet_1_0__leaf_net504),
    .A1(net496),
    .A2(clknet_1_0__leaf_net503),
    .A3(net371),
    .S0(net498),
    .S1(net850),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(clknet_1_0__leaf_net503),
    .A1(net494),
    .A2(net498),
    .A3(net480),
    .S0(net848),
    .S1(net850),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c682 (.A0(clknet_1_1__leaf_net488),
    .A1(clknet_1_0__leaf_net391),
    .A2(net252),
    .A3(net1127),
    .S0(net1126),
    .S1(net847),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c683 (.A0(net894),
    .A1(clknet_1_0__leaf_net261),
    .A2(net1062),
    .A3(net1055),
    .S0(net700),
    .S1(clknet_1_1__leaf_net743),
    .X(net508));
 sky130_fd_sc_hd__mux4_1 c684 (.A0(net1060),
    .A1(net1073),
    .A2(net500),
    .A3(net652),
    .S0(net753),
    .S1(net825),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c685 (.A0(net376),
    .A1(clknet_1_1__leaf_net503),
    .A2(net499),
    .A3(net1063),
    .S0(clknet_1_1__leaf_net704),
    .S1(clknet_1_1__leaf_net743),
    .X(net510));
 sky130_fd_sc_hd__mux4_2 c686 (.A0(net1117),
    .A1(net1120),
    .A2(net1115),
    .A3(net264),
    .S0(net789),
    .S1(net851),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c687 (.A0(net499),
    .A1(clknet_1_1__leaf_net503),
    .A2(net397),
    .A3(net786),
    .S0(net829),
    .S1(net853),
    .X(net512));
 sky130_fd_sc_hd__mux4_1 c688 (.A0(net1103),
    .A1(net1121),
    .A2(net894),
    .A3(clknet_1_0__leaf_net503),
    .S0(net874),
    .S1(net753),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c689 (.A0(clknet_1_0__leaf_net503),
    .A1(net397),
    .A2(net1120),
    .A3(net498),
    .S0(net1110),
    .S1(net847),
    .X(net514));
 sky130_fd_sc_hd__mux4_1 c690 (.A0(net1069),
    .A1(net1052),
    .A2(net59),
    .A3(net39),
    .S0(net1170),
    .S1(net1139),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c691 (.A0(clknet_1_0__leaf_net513),
    .A1(net1117),
    .A2(net1100),
    .A3(net652),
    .S0(net813),
    .S1(clknet_1_0__leaf_net820),
    .X(net516));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(net500),
    .A1(net53),
    .A2(net869),
    .A3(net367),
    .S0(net609),
    .S1(net789),
    .X(net517));
 sky130_fd_sc_hd__mux4_1 c693 (.A0(net380),
    .A1(net397),
    .A2(clknet_1_0__leaf_net261),
    .A3(net1121),
    .S0(net849),
    .S1(net856),
    .X(net518));
 sky130_fd_sc_hd__mux4_1 c694 (.A0(net482),
    .A1(net1097),
    .A2(net1115),
    .A3(clknet_1_0__leaf_net513),
    .S0(net1119),
    .S1(net855),
    .X(net519));
 sky130_fd_sc_hd__mux4_1 c695 (.A0(clknet_1_1__leaf_net398),
    .A1(clknet_1_1__leaf_net513),
    .A2(net1126),
    .A3(net594),
    .S0(net847),
    .S1(net856),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 c696 (.A0(clknet_1_0__leaf_net516),
    .A1(clknet_1_1__leaf_net393),
    .A2(net894),
    .A3(net500),
    .S0(net786),
    .S1(net856),
    .X(net521));
 sky130_fd_sc_hd__mux4_1 c697 (.A0(clknet_1_0__leaf_net390),
    .A1(net1126),
    .A2(net500),
    .A3(net1061),
    .S0(net669),
    .S1(net856),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(net494),
    .A1(clknet_1_1__leaf_net503),
    .A2(net675),
    .A3(clknet_1_1__leaf_net820),
    .S0(net852),
    .S1(net856),
    .X(net523));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(clknet_1_1__leaf_net398),
    .A1(net1061),
    .A2(net614),
    .A3(net675),
    .S0(net691),
    .S1(net780),
    .X(net524));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(clknet_1_1__leaf_net513),
    .A1(net251),
    .A2(net511),
    .A3(net706),
    .S0(net753),
    .S1(net856),
    .X(net525));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(clknet_1_1__leaf_net503),
    .A1(clknet_1_0__leaf_net525),
    .A2(net669),
    .A3(net673),
    .S0(net847),
    .S1(net848),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(clknet_1_1__leaf_net525),
    .A1(net499),
    .A2(net368),
    .A3(net1108),
    .S0(net1110),
    .S1(net626),
    .X(net527));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(net520),
    .A1(net1120),
    .A2(net511),
    .A3(net1063),
    .S0(net595),
    .S1(net691),
    .X(net528));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net510),
    .A1(net1127),
    .A2(net264),
    .A3(net1116),
    .S0(clknet_1_1__leaf_net820),
    .S1(net1084),
    .X(net529));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(clknet_1_0__leaf_net391),
    .A1(clknet_1_0__leaf_net431),
    .A2(net53),
    .A3(net491),
    .S0(net829),
    .S1(net837),
    .X(net530));
 sky130_fd_sc_hd__mux4_1 c706 (.A0(clknet_1_0__leaf_net506),
    .A1(net1119),
    .A2(net55),
    .A3(net920),
    .S0(net885),
    .S1(net908),
    .X(net531));
 sky130_fd_sc_hd__mux4_1 c707 (.A0(net303),
    .A1(net905),
    .A2(net1065),
    .A3(net187),
    .S0(net625),
    .S1(net1084),
    .X(net532));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(clknet_1_0__leaf_net529),
    .A1(net424),
    .A2(net780),
    .A3(net796),
    .S0(net837),
    .S1(net857),
    .X(net533));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(net495),
    .A1(net894),
    .A2(net905),
    .A3(clknet_1_1__leaf_net523),
    .S0(net856),
    .S1(clknet_1_0__leaf_net859),
    .X(net534));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net1065),
    .A1(net903),
    .A2(net609),
    .A3(net780),
    .S0(clknet_1_1__leaf_net800),
    .S1(net826),
    .X(net535));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net905),
    .A1(net46),
    .A2(net1059),
    .A3(net715),
    .S0(net837),
    .S1(net857),
    .X(net536));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(clknet_1_0__leaf_net523),
    .A1(clknet_1_1__leaf_net506),
    .A2(net53),
    .A3(net792),
    .S0(net797),
    .S1(net848),
    .X(net537));
 sky130_fd_sc_hd__mux4_1 c713 (.A0(clknet_1_0__leaf_net430),
    .A1(net974),
    .A2(net1062),
    .A3(net814),
    .S0(clknet_1_0__leaf_net838),
    .S1(clknet_1_0__leaf_net860),
    .X(net538));
 sky130_fd_sc_hd__mux4_2 c714 (.A0(net368),
    .A1(net908),
    .A2(net495),
    .A3(net285),
    .S0(net1172),
    .S1(net691),
    .X(net977));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net491),
    .A1(net412),
    .A2(net837),
    .A3(clknet_1_0__leaf_net839),
    .S0(net857),
    .S1(clknet_1_0__leaf_net860),
    .X(net539));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net1172),
    .A1(net905),
    .A2(net977),
    .A3(net1063),
    .S0(net367),
    .S1(net490),
    .X(net540));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net1073),
    .A1(net920),
    .A2(clknet_1_1__leaf_net277),
    .A3(clknet_1_1__leaf_net291),
    .S0(net798),
    .S1(clknet_1_1__leaf_net859),
    .X(net541));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(clknet_1_0__leaf_net539),
    .A1(clknet_1_0__leaf_net430),
    .A2(net825),
    .A3(net848),
    .S0(net853),
    .S1(net857),
    .X(net542));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net478),
    .A1(clknet_1_0__leaf_net539),
    .A2(net1116),
    .A3(net874),
    .S0(net785),
    .S1(net837),
    .X(net543));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net534),
    .A1(net538),
    .A2(net977),
    .A3(clknet_1_1__leaf_net430),
    .S0(clknet_1_1__leaf_net539),
    .S1(net1059),
    .X(net544));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net880),
    .A1(clknet_1_1__leaf_net391),
    .A2(net877),
    .A3(net1101),
    .S0(net973),
    .S1(clknet_1_0__leaf_net859),
    .X(net545));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net543),
    .A1(net59),
    .A2(net315),
    .A3(net877),
    .S0(net673),
    .S1(clknet_1_1__leaf_net858),
    .X(net546));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(clknet_1_1__leaf_net277),
    .A1(clknet_1_1__leaf_net539),
    .A2(net494),
    .A3(net1061),
    .S0(net857),
    .S1(clknet_1_1__leaf_net858),
    .X(net547));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(clknet_1_1__leaf_net529),
    .A1(net1053),
    .A2(net668),
    .A3(net833),
    .S0(clknet_1_1__leaf_net858),
    .S1(clknet_1_0__leaf_net860),
    .X(net548));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net188),
    .A1(clknet_1_0__leaf_net529),
    .A2(net397),
    .A3(net673),
    .S0(net762),
    .S1(clknet_1_0__leaf_net860),
    .X(net549));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net303),
    .A1(net949),
    .A2(net648),
    .A3(net1083),
    .S0(net780),
    .S1(net829),
    .X(net550));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(clknet_1_1__leaf_net215),
    .A1(net511),
    .A2(net903),
    .A3(net772),
    .S0(clknet_1_1__leaf_net818),
    .S1(net863),
    .X(net551));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net1069),
    .A1(net265),
    .A2(clknet_1_1__leaf_net393),
    .A3(net1083),
    .S0(net762),
    .S1(net1084),
    .X(net1030));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(clknet_1_1__leaf_net519),
    .A1(clknet_1_1__leaf_net261),
    .A2(net1087),
    .A3(net1105),
    .S0(net649),
    .S1(clknet_1_1__leaf_net838),
    .X(net552));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net908),
    .A1(clknet_1_1__leaf_net328),
    .A2(net265),
    .A3(net747),
    .S0(clknet_1_1__leaf_net818),
    .S1(net861),
    .X(net553));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net941),
    .A1(clknet_1_0__leaf_net324),
    .A2(clknet_1_1__leaf_net635),
    .A3(net721),
    .S0(clknet_1_0__leaf_net858),
    .S1(clknet_1_1__leaf_net860),
    .X(net554));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(clknet_1_0__leaf_net456),
    .A1(net971),
    .A2(clknet_1_1__leaf_net328),
    .A3(net772),
    .S0(net789),
    .S1(clknet_1_0__leaf_net858),
    .X(net555));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net412),
    .A1(net941),
    .A2(net903),
    .A3(clknet_1_1__leaf_net1022),
    .S0(net684),
    .S1(clknet_1_1__leaf_net704),
    .X(net556));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(net894),
    .A1(net55),
    .A2(net1059),
    .A3(clknet_1_1__leaf_net860),
    .S0(net862),
    .S1(net865),
    .X(net557));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net78),
    .A1(net690),
    .A2(net829),
    .A3(net851),
    .S0(net864),
    .S1(net866),
    .X(net558));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(clknet_1_1__leaf_net504),
    .A1(net1119),
    .A2(net941),
    .A3(net558),
    .S0(clknet_1_1__leaf_net818),
    .S1(net856),
    .X(net559));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(clknet_1_0__leaf_net393),
    .A1(clknet_1_0__leaf_net505),
    .A2(net629),
    .A3(net674),
    .S0(clknet_1_1__leaf_net743),
    .S1(net863),
    .X(net560));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net252),
    .A1(net326),
    .A2(net673),
    .A3(net728),
    .S0(net1084),
    .S1(net857),
    .X(net561));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(clknet_1_1__leaf_net435),
    .A1(clknet_1_1__leaf_net516),
    .A2(net265),
    .A3(net674),
    .S0(clknet_1_1__leaf_net743),
    .S1(net747),
    .X(net562));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(net556),
    .A1(net558),
    .A2(clknet_1_1__leaf_net456),
    .A3(net412),
    .S0(net808),
    .S1(net994),
    .X(net563));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(net542),
    .A1(net412),
    .A2(net65),
    .A3(net40),
    .S0(net684),
    .S1(net772),
    .X(net564));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(clknet_1_0__leaf_net564),
    .A1(net941),
    .A2(net686),
    .A3(net762),
    .S0(net854),
    .S1(clknet_1_1__leaf_net859),
    .X(net565));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(clknet_1_0__leaf_net519),
    .A1(clknet_1_0__leaf_net564),
    .A2(net1069),
    .A3(clknet_1_1__leaf_net635),
    .S0(net686),
    .S1(net805),
    .X(net566));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(clknet_1_1__leaf_net505),
    .A1(clknet_1_1__leaf_net564),
    .A2(net1063),
    .A3(net692),
    .S0(clknet_1_1__leaf_net860),
    .S1(net862),
    .X(net567));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(clknet_1_1__leaf_net564),
    .A1(net686),
    .A2(net707),
    .A3(clknet_1_1__leaf_net818),
    .S0(net1084),
    .S1(net864),
    .X(net568));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net326),
    .A1(clknet_1_1__leaf_net564),
    .A2(net684),
    .A3(net685),
    .S0(net973),
    .S1(net692),
    .X(net569));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(net326),
    .A1(clknet_1_1__leaf_net324),
    .A2(net1061),
    .A3(net690),
    .S0(clknet_1_1__leaf_net743),
    .S1(clknet_1_1__leaf_net860),
    .X(net570));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net899),
    .A1(net1063),
    .A2(clknet_1_1__leaf_net681),
    .A3(net712),
    .S0(net811),
    .S1(net845),
    .X(net571));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net1101),
    .A1(net1097),
    .A2(net961),
    .A3(net668),
    .S0(net693),
    .S1(net811),
    .X(net572));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(clknet_1_1__leaf_net390),
    .A1(net59),
    .A2(net1059),
    .A3(clknet_1_1__leaf_net241),
    .S0(net1079),
    .S1(net868),
    .X(net573));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net252),
    .A1(net1065),
    .A2(net908),
    .A3(net902),
    .S0(net1105),
    .S1(net827),
    .X(net574));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net65),
    .A1(net143),
    .A2(clknet_1_1__leaf_net464),
    .A3(net973),
    .S0(net689),
    .S1(net693),
    .X(net575));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(clknet_1_0__leaf_net241),
    .A1(net572),
    .A2(clknet_1_1__leaf_net390),
    .A3(net920),
    .S0(net747),
    .S1(net826),
    .X(net576));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net285),
    .A1(net1059),
    .A2(net679),
    .A3(net857),
    .S0(net867),
    .S1(net868),
    .X(net577));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net26),
    .A1(net891),
    .A2(net877),
    .A3(net797),
    .S0(clknet_1_0__leaf_net801),
    .S1(net852),
    .X(net578));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net877),
    .A1(net961),
    .A2(clknet_1_0__leaf_net969),
    .A3(net712),
    .S0(net772),
    .S1(net867),
    .X(net579));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net535),
    .A1(clknet_1_1__leaf_net100),
    .A2(net892),
    .A3(net690),
    .S0(clknet_1_1__leaf_net704),
    .S1(net857),
    .X(net580));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(clknet_1_1__leaf_net328),
    .A1(net903),
    .A2(net476),
    .A3(net1070),
    .S0(net40),
    .S1(net674),
    .X(net581));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net908),
    .A1(clknet_1_1__leaf_net458),
    .A2(net874),
    .A3(net687),
    .S0(net762),
    .S1(clknet_1_1__leaf_net840),
    .X(net582));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net874),
    .A1(net40),
    .A2(net578),
    .A3(clknet_1_1__leaf_net458),
    .S0(net1065),
    .S1(net675),
    .X(net583));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(clknet_1_1__leaf_net261),
    .A1(net1103),
    .A2(net580),
    .A3(net26),
    .S0(net674),
    .S1(net685),
    .X(net584));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(clknet_1_1__leaf_net100),
    .A1(net1105),
    .A2(net554),
    .A3(net59),
    .S0(net687),
    .S1(clknet_1_0__leaf_net839),
    .X(net585));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(net315),
    .A1(net78),
    .A2(net1098),
    .A3(clknet_1_1__leaf_net681),
    .S0(net808),
    .S1(net811),
    .X(net586));
 sky130_fd_sc_hd__mux4_1 c764 (.A0(net377),
    .A1(net913),
    .A2(net762),
    .A3(clknet_1_1__leaf_net801),
    .S0(clknet_1_1__leaf_net840),
    .S1(net854),
    .X(net587));
 sky130_fd_sc_hd__mux4_1 c765 (.A0(net265),
    .A1(clknet_1_1__leaf_net324),
    .A2(net688),
    .A3(net690),
    .S0(net721),
    .S1(net856),
    .X(net588));
 sky130_fd_sc_hd__mux4_1 c766 (.A0(net949),
    .A1(net571),
    .A2(net680),
    .A3(net684),
    .S0(net685),
    .S1(net1079),
    .X(net589));
 sky130_fd_sc_hd__mux4_1 c767 (.A0(net588),
    .A1(net574),
    .A2(clknet_1_0__leaf_net681),
    .A3(net686),
    .S0(net773),
    .S1(net856),
    .X(net590));
 sky130_fd_sc_hd__mux4_1 c768 (.A0(net589),
    .A1(clknet_1_1__leaf_net460),
    .A2(net902),
    .A3(net587),
    .S0(net1040),
    .S1(net680),
    .X(net591));
 sky130_fd_sc_hd__mux4_1 c769 (.A0(clknet_1_1__leaf_net291),
    .A1(net46),
    .A2(net629),
    .A3(net675),
    .S0(clknet_1_0__leaf_net681),
    .S1(net685),
    .X(net592));
 sky130_fd_sc_hd__xnor2_1 merge790 (.A(net457),
    .B(net459),
    .Y(net593));
 sky130_fd_sc_hd__dfrbp_1 merge791 (.CLK(clknet_leaf_13_clk),
    .D(net508),
    .RESET_B(net515),
    .Q(net595),
    .Q_N(net594));
 sky130_fd_sc_hd__xnor2_1 merge792 (.A(net226),
    .B(net207),
    .Y(net596));
 sky130_fd_sc_hd__dfrbp_2 merge793 (.CLK(clknet_leaf_40_clk),
    .D(net101),
    .RESET_B(net89),
    .Q(net997),
    .Q_N(net597));
 sky130_fd_sc_hd__dfrtn_1 merge794 (.CLK_N(clknet_leaf_46_clk),
    .D(net63),
    .RESET_B(net51),
    .Q(net598));
 sky130_fd_sc_hd__xnor2_1 merge795 (.A(net550),
    .B(net551),
    .Y(net599));
 sky130_fd_sc_hd__dfrtp_4 merge796 (.CLK(clknet_leaf_9_clk),
    .D(net378),
    .RESET_B(net369),
    .Q(net600));
 sky130_fd_sc_hd__xnor2_1 merge797 (.A(net395),
    .B(net402),
    .Y(net601));
 sky130_fd_sc_hd__xnor2_1 merge798 (.A(net355),
    .B(net356),
    .Y(net602));
 sky130_fd_sc_hd__xnor2_1 merge799 (.A(net437),
    .B(net440),
    .Y(net603));
 sky130_fd_sc_hd__xnor2_1 merge800 (.A(net204),
    .B(net205),
    .Y(net604));
 sky130_fd_sc_hd__dfrtp_4 merge801 (.CLK(clknet_leaf_2_clk),
    .D(net175),
    .RESET_B(net182),
    .Q(net605));
 sky130_fd_sc_hd__xnor2_1 merge802 (.A(net327),
    .B(net334),
    .Y(net606));
 sky130_fd_sc_hd__xnor2_1 merge803 (.A(net227),
    .B(net235),
    .Y(net607));
 sky130_fd_sc_hd__dfrtp_4 merge804 (.CLK(clknet_leaf_36_clk),
    .D(net4),
    .RESET_B(net6),
    .Q(net1023));
 sky130_fd_sc_hd__dfsbp_2 merge805 (.CLK(clknet_leaf_11_clk),
    .SET_B(net479),
    .Q(net609),
    .Q_N(net483));
 sky130_fd_sc_hd__dfsbp_2 merge806 (.CLK(clknet_leaf_48_clk),
    .D(net30),
    .SET_B(net32),
    .Q(net611),
    .Q_N(net610));
 sky130_fd_sc_hd__dfstp_1 merge807 (.CLK(clknet_leaf_45_clk),
    .SET_B(net79),
    .Q(net87));
 sky130_fd_sc_hd__xnor2_1 merge808 (.A(net127),
    .B(net129),
    .Y(net613));
 sky130_fd_sc_hd__dfstp_2 merge809 (.CLK(clknet_leaf_3_clk),
    .D(net300),
    .SET_B(net283),
    .Q(net614));
 sky130_fd_sc_hd__xnor2_1 merge810 (.A(net531),
    .B(net532),
    .Y(net615));
 sky130_fd_sc_hd__dfstp_2 merge811 (.CLK(clknet_leaf_7_clk),
    .D(net275),
    .SET_B(net250),
    .Q(net616));
 sky130_fd_sc_hd__dlrbn_2 merge812 (.D(net158),
    .GATE_N(clknet_leaf_1_clk),
    .RESET_B(net139),
    .Q(net618),
    .Q_N(net617));
 sky130_fd_sc_hd__dlrbn_1 merge813 (.D(net119),
    .GATE_N(clknet_leaf_35_clk),
    .RESET_B(net126),
    .Q(net619),
    .Q_N(net984));
 sky130_fd_sc_hd__xnor2_1 merge814 (.A(net592),
    .B(net573),
    .Y(net620));
 sky130_fd_sc_hd__dlrbp_1 merge815 (.D(net309),
    .GATE(clknet_leaf_4_clk),
    .RESET_B(net313),
    .Q(net622),
    .Q_N(net621));
 sky130_fd_sc_hd__xnor2_1 merge816 (.A(net21),
    .B(net10),
    .Y(net623));
 sky130_fd_sc_hd__xnor2_1 merge817 (.A(net434),
    .B(net415),
    .Y(net624));
 sky130_fd_sc_hd__dlrbp_1 merge818 (.D(net526),
    .GATE(clknet_leaf_14_clk),
    .RESET_B(net524),
    .Q(net626),
    .Q_N(net625));
 sky130_fd_sc_hd__dlrtn_4 merge819 (.D(net160),
    .GATE_N(clknet_leaf_2_clk),
    .RESET_B(net168),
    .Q(net627));
 sky130_fd_sc_hd__dlrtn_2 merge820 (.D(net109),
    .GATE_N(clknet_leaf_37_clk),
    .RESET_B(net107),
    .Q(net1004));
 sky130_fd_sc_hd__xnor2_1 merge821 (.A(net522),
    .B(net521),
    .Y(net628));
 sky130_fd_sc_hd__dlrtn_1 merge822 (.D(net64),
    .GATE_N(clknet_leaf_46_clk),
    .Q(net66));
 sky130_fd_sc_hd__xnor2_1 merge823 (.A(net236),
    .B(net243),
    .Y(net630));
 sky130_fd_sc_hd__dlrtp_1 merge824 (.D(net209),
    .GATE(clknet_leaf_39_clk),
    .RESET_B(net216),
    .Q(net631));
 sky130_fd_sc_hd__xnor2_1 merge825 (.A(net359),
    .B(net449),
    .Y(net632));
 sky130_fd_sc_hd__dlrtp_1 merge826 (.D(net131),
    .GATE(clknet_leaf_36_clk),
    .RESET_B(net18),
    .Q(net1046));
 sky130_fd_sc_hd__dlrtp_1 merge827 (.D(net11),
    .GATE(clknet_leaf_36_clk),
    .RESET_B(net613),
    .Q(net1047));
 sky130_fd_sc_hd__edfxbp_1 merge828 (.CLK(clknet_leaf_34_clk),
    .D(net110),
    .DE(net124),
    .Q(net1033),
    .Q_N(net633));
 sky130_fd_sc_hd__edfxtp_1 merge829 (.CLK(clknet_leaf_17_clk),
    .D(net429),
    .DE(net418),
    .Q(net634));
 sky130_fd_sc_hd__sdlclkp_1 merge830 (.CLK(clknet_leaf_45_clk),
    .GATE(net85),
    .SCE(net81),
    .GCLK(net635));
 sky130_fd_sc_hd__sdlclkp_2 merge831 (.CLK(clknet_leaf_25_clk),
    .GATE(net472),
    .SCE(net471),
    .GCLK(net970));
 sky130_fd_sc_hd__xnor2_1 merge832 (.A(net239),
    .B(net17),
    .Y(net636));
 sky130_fd_sc_hd__sdlclkp_4 merge833 (.CLK(clknet_leaf_31_clk),
    .GATE(net607),
    .SCE(net632),
    .GCLK(net637));
 sky130_fd_sc_hd__xnor2_1 merge834 (.A(net544),
    .B(net570),
    .Y(net638));
 sky130_fd_sc_hd__xnor2_1 merge835 (.A(net536),
    .B(net591),
    .Y(net639));
 sky130_fd_sc_hd__dfrbp_1 merge836 (.CLK(clknet_leaf_31_clk),
    .D(net347),
    .RESET_B(net338),
    .Q(net641),
    .Q_N(net640));
 sky130_fd_sc_hd__xnor2_1 merge837 (.A(net620),
    .B(net454),
    .Y(net642));
 sky130_fd_sc_hd__xnor2_1 merge838 (.A(net467),
    .B(net590),
    .Y(net643));
 sky130_fd_sc_hd__xnor2_1 merge839 (.A(net443),
    .B(net466),
    .Y(net644));
 sky130_fd_sc_hd__xnor2_1 merge840 (.A(net565),
    .B(net586),
    .Y(net645));
 sky130_fd_sc_hd__xnor2_1 merge841 (.A(net549),
    .B(net548),
    .Y(net646));
 sky130_fd_sc_hd__xnor2_1 merge842 (.A(net540),
    .B(net569),
    .Y(net647));
 sky130_fd_sc_hd__dfrbp_1 merge843 (.CLK(clknet_leaf_21_clk),
    .D(net545),
    .RESET_B(net541),
    .Q(net649),
    .Q_N(net648));
 sky130_fd_sc_hd__xnor2_1 merge844 (.A(net455),
    .B(net446),
    .Y(net650));
 sky130_fd_sc_hd__dfrtn_1 merge845 (.CLK_N(clknet_leaf_16_clk),
    .RESET_B(net407),
    .Q(net651));
 sky130_fd_sc_hd__dfrtp_1 merge846 (.CLK(clknet_leaf_4_clk),
    .RESET_B(net295),
    .Q(net302));
 sky130_fd_sc_hd__dfrtp_4 merge847 (.CLK(clknet_leaf_42_clk),
    .D(net203),
    .RESET_B(net196),
    .Q(net1014));
 sky130_fd_sc_hd__xnor2_1 merge848 (.A(net575),
    .B(net576),
    .Y(net653));
 sky130_fd_sc_hd__xnor2_1 merge849 (.A(net321),
    .B(net602),
    .Y(net654));
 sky130_fd_sc_hd__dfrtp_1 merge850 (.CLK(clknet_leaf_36_clk),
    .D(net16),
    .RESET_B(net15),
    .Q(net1045));
 sky130_fd_sc_hd__dfsbp_1 merge851 (.CLK(clknet_leaf_18_clk),
    .SET_B(net320),
    .Q(net656),
    .Q_N(net322));
 sky130_fd_sc_hd__xnor2_1 merge852 (.A(net553),
    .B(net585),
    .Y(net657));
 sky130_fd_sc_hd__dfsbp_2 merge853 (.CLK(clknet_leaf_30_clk),
    .D(net342),
    .SET_B(net606),
    .Q(net1012),
    .Q_N(net658));
 sky130_fd_sc_hd__xnor2_1 merge854 (.A(net566),
    .B(net584),
    .Y(net659));
 sky130_fd_sc_hd__dfstp_2 merge855 (.CLK(clknet_leaf_24_clk),
    .D(net444),
    .SET_B(net643),
    .Q(net1040));
 sky130_fd_sc_hd__dfstp_1 merge856 (.CLK(clknet_leaf_27_clk),
    .D(net445),
    .SET_B(net650),
    .Q(net660));
 sky130_fd_sc_hd__dfstp_1 merge857 (.CLK(clknet_leaf_32_clk),
    .D(net366),
    .SET_B(net630),
    .Q(net661));
 sky130_fd_sc_hd__dlrbn_1 merge858 (.D(net333),
    .GATE_N(clknet_leaf_26_clk),
    .RESET_B(net344),
    .Q(net663),
    .Q_N(net662));
 sky130_fd_sc_hd__dlrbn_1 merge859 (.D(net354),
    .GATE_N(clknet_leaf_32_clk),
    .RESET_B(net351),
    .Q(net665),
    .Q_N(net664));
 sky130_fd_sc_hd__xnor2_1 merge860 (.A(net582),
    .B(net567),
    .Y(net666));
 sky130_fd_sc_hd__xnor2_1 merge861 (.A(net581),
    .B(net568),
    .Y(net667));
 sky130_fd_sc_hd__dlrbp_1 merge862 (.D(net518),
    .GATE(clknet_leaf_13_clk),
    .RESET_B(net647),
    .Q(net669),
    .Q_N(net668));
 sky130_fd_sc_hd__xnor2_1 merge863 (.A(net583),
    .B(net577),
    .Y(net670));
 sky130_fd_sc_hd__dlrbp_1 merge864 (.D(net234),
    .GATE(clknet_leaf_30_clk),
    .RESET_B(net210),
    .Q(net672),
    .Q_N(net671));
 sky130_fd_sc_hd__dlrtn_1 merge865 (.D(net512),
    .GATE_N(clknet_leaf_14_clk),
    .RESET_B(net646),
    .Q(net673));
 sky130_fd_sc_hd__dlrtn_1 merge866 (.D(net670),
    .GATE_N(clknet_leaf_20_clk),
    .RESET_B(net552),
    .Q(net674));
 sky130_fd_sc_hd__dlrtn_1 merge867 (.D(net644),
    .GATE_N(clknet_leaf_27_clk),
    .RESET_B(net593),
    .Q(net993));
 sky130_fd_sc_hd__dlrtp_1 merge868 (.D(net639),
    .GATE(clknet_leaf_21_clk),
    .RESET_B(net628),
    .Q(net675));
 sky130_fd_sc_hd__dlrtp_2 merge869 (.D(net230),
    .GATE(clknet_leaf_37_clk),
    .RESET_B(net219),
    .Q(net676));
 sky130_fd_sc_hd__dlrtp_1 merge870 (.D(net603),
    .GATE(clknet_leaf_28_clk),
    .RESET_B(net441),
    .Q(net677));
 sky130_fd_sc_hd__edfxbp_1 merge871 (.CLK(clknet_leaf_27_clk),
    .D(net463),
    .DE(net450),
    .Q(net679),
    .Q_N(net678));
 sky130_fd_sc_hd__edfxtp_1 merge872 (.CLK(clknet_leaf_24_clk),
    .D(net452),
    .DE(net645),
    .Q(net680));
 sky130_fd_sc_hd__sdlclkp_1 merge873 (.CLK(clknet_leaf_30_clk),
    .GATE(net596),
    .SCE(net222),
    .GCLK(net1022));
 sky130_fd_sc_hd__sdlclkp_2 merge874 (.CLK(clknet_leaf_7_clk),
    .GATE(net276),
    .SCE(net654),
    .GCLK(net999));
 sky130_fd_sc_hd__sdlclkp_4 merge875 (.CLK(clknet_leaf_20_clk),
    .GATE(net599),
    .SCE(net659),
    .GCLK(net681));
 sky130_fd_sc_hd__dfrbp_2 merge876 (.CLK(clknet_leaf_35_clk),
    .D(net121),
    .RESET_B(net130),
    .Q(net682),
    .Q_N(net1018));
 sky130_fd_sc_hd__dfrbp_2 merge877 (.CLK(clknet_leaf_36_clk),
    .D(net123),
    .RESET_B(net623),
    .Q(net683),
    .Q_N(net1031));
 sky130_fd_sc_hd__dfrtn_1 merge878 (.CLK_N(clknet_leaf_23_clk),
    .D(net453),
    .RESET_B(net657),
    .Q(net684));
 sky130_fd_sc_hd__dfrtp_2 merge879 (.CLK(clknet_leaf_22_clk),
    .D(net561),
    .RESET_B(net667),
    .Q(net685));
 sky130_fd_sc_hd__dfrtp_2 merge880 (.CLK(clknet_leaf_23_clk),
    .D(net563),
    .RESET_B(net666),
    .Q(net686));
 sky130_fd_sc_hd__dfrtp_4 merge881 (.CLK(clknet_leaf_22_clk),
    .D(net638),
    .RESET_B(net562),
    .Q(net973));
 sky130_fd_sc_hd__dfsbp_1 merge882 (.CLK(clknet_leaf_19_clk),
    .D(net451),
    .SET_B(net653),
    .Q(net980),
    .Q_N(net687));
 sky130_fd_sc_hd__dfsbp_1 merge883 (.CLK(clknet_leaf_24_clk),
    .D(net475),
    .SET_B(net642),
    .Q(net689),
    .Q_N(net688));
 sky130_fd_sc_hd__dfstp_2 merge884 (.CLK(clknet_leaf_35_clk),
    .D(net238),
    .SET_B(net1152),
    .Q(net1036));
 sky130_fd_sc_hd__dfstp_1 merge885 (.CLK(clknet_leaf_23_clk),
    .D(net527),
    .SET_B(net579),
    .Q(net690));
 sky130_fd_sc_hd__dfstp_4 merge886 (.CLK(clknet_leaf_42_clk),
    .D(net604),
    .SET_B(net176),
    .Q(net691));
 sky130_fd_sc_hd__dlrbn_1 merge887 (.D(net615),
    .GATE_N(clknet_leaf_22_clk),
    .RESET_B(net559),
    .Q(net693),
    .Q_N(net692));
 sky130_fd_sc_hd__dlrbn_1 merge888 (.D(net636),
    .GATE_N(clknet_leaf_32_clk),
    .RESET_B(net246),
    .Q(net988),
    .Q_N(net694));
 sky130_fd_sc_hd__dlrbp_1 merge889 (.D(net601),
    .GATE(clknet_leaf_17_clk),
    .RESET_B(net624),
    .Q(net695),
    .Q_N(net982));
 sky130_fd_sc_hd__dlxtp_1 s1000 (.D(net414),
    .GATE(clknet_2_1__leaf_clk),
    .Q(net830));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s1001 (.D(net417),
    .SLEEP_B(clknet_leaf_18_clk),
    .Q(net831));
 sky130_fd_sc_hd__dfxbp_1 s1002 (.CLK(clknet_leaf_17_clk),
    .D(net419),
    .Q(net833),
    .Q_N(net832));
 sky130_fd_sc_hd__dfxbp_1 s1003 (.CLK(clknet_leaf_17_clk),
    .D(net420),
    .Q(net835),
    .Q_N(net834));
 sky130_fd_sc_hd__dfxtp_1 s1004 (.CLK(clknet_leaf_17_clk),
    .D(net421),
    .Q(net836));
 sky130_fd_sc_hd__dfxtp_2 s1005 (.CLK(clknet_leaf_19_clk),
    .D(net423),
    .Q(net837));
 sky130_fd_sc_hd__dfxtp_2 s1006 (.CLK(clknet_leaf_14_clk),
    .D(net426),
    .Q(net989));
 sky130_fd_sc_hd__dlclkp_1 s1007 (.CLK(clknet_leaf_19_clk),
    .GATE(net427),
    .GCLK(net838));
 sky130_fd_sc_hd__dlclkp_2 s1008 (.CLK(clknet_leaf_17_clk),
    .GATE(net428),
    .GCLK(net839));
 sky130_fd_sc_hd__dlclkp_4 s1009 (.CLK(clknet_leaf_26_clk),
    .GATE(net438),
    .GCLK(net840));
 sky130_fd_sc_hd__dlxbn_1 s1010 (.D(net447),
    .GATE_N(clknet_leaf_27_clk),
    .Q(net842),
    .Q_N(net841));
 sky130_fd_sc_hd__dlxbn_2 s1011 (.D(net448),
    .GATE_N(clknet_leaf_24_clk),
    .Q(net994),
    .Q_N(net843));
 sky130_fd_sc_hd__dlxbp_1 s1012 (.D(net461),
    .GATE(clknet_leaf_26_clk),
    .Q(net845),
    .Q_N(net844));
 sky130_fd_sc_hd__dlxtn_1 s1013 (.D(net469),
    .GATE_N(clknet_leaf_25_clk),
    .Q(net846));
 sky130_fd_sc_hd__dlxtn_2 s1014 (.D(net489),
    .GATE_N(clknet_leaf_11_clk),
    .Q(net847));
 sky130_fd_sc_hd__dlxtn_2 s1015 (.D(net492),
    .GATE_N(clknet_leaf_12_clk),
    .Q(net848));
 sky130_fd_sc_hd__dlxtp_1 s1016 (.D(net501),
    .GATE(clknet_leaf_12_clk),
    .Q(net849));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s1017 (.D(net502),
    .SLEEP_B(clknet_leaf_12_clk),
    .Q(net850));
 sky130_fd_sc_hd__dfxbp_1 s1018 (.CLK(clknet_leaf_13_clk),
    .D(net507),
    .Q(net852),
    .Q_N(net851));
 sky130_fd_sc_hd__dfxbp_1 s1019 (.CLK(clknet_leaf_15_clk),
    .D(net509),
    .Q(net854),
    .Q_N(net853));
 sky130_fd_sc_hd__dfxtp_1 s1020 (.CLK(clknet_leaf_12_clk),
    .D(net514),
    .Q(net855));
 sky130_fd_sc_hd__dfxtp_4 s1021 (.CLK(clknet_leaf_13_clk),
    .D(net517),
    .Q(net856));
 sky130_fd_sc_hd__dfxtp_4 s1022 (.CLK(clknet_leaf_14_clk),
    .D(net528),
    .Q(net857));
 sky130_fd_sc_hd__dlclkp_1 s1023 (.CLK(clknet_leaf_21_clk),
    .GATE(net530),
    .GCLK(net858));
 sky130_fd_sc_hd__dlclkp_2 s1024 (.CLK(clknet_leaf_15_clk),
    .GATE(net533),
    .GCLK(net859));
 sky130_fd_sc_hd__dlclkp_4 s1025 (.CLK(clknet_leaf_14_clk),
    .GATE(net537),
    .GCLK(net860));
 sky130_fd_sc_hd__dlxbn_1 s1026 (.D(net546),
    .GATE_N(clknet_leaf_22_clk),
    .Q(net862),
    .Q_N(net861));
 sky130_fd_sc_hd__dlxbn_1 s1027 (.D(net547),
    .GATE_N(clknet_leaf_21_clk),
    .Q(net864),
    .Q_N(net863));
 sky130_fd_sc_hd__dlxbp_1 s1028 (.D(net555),
    .GATE(clknet_leaf_22_clk),
    .Q(net866),
    .Q_N(net865));
 sky130_fd_sc_hd__dlxtn_1 s1029 (.D(net557),
    .GATE_N(clknet_leaf_23_clk),
    .Q(net867));
 sky130_fd_sc_hd__dlxtn_1 s1030 (.D(net560),
    .GATE_N(clknet_leaf_23_clk),
    .Q(net868));
 sky130_fd_sc_hd__dfxbp_2 s890 (.CLK(clknet_leaf_48_clk),
    .D(net31),
    .Q(net697),
    .Q_N(net696));
 sky130_fd_sc_hd__dfxbp_2 s891 (.CLK(clknet_leaf_49_clk),
    .D(net33),
    .Q(net699),
    .Q_N(net698));
 sky130_fd_sc_hd__dfxtp_4 s892 (.CLK(clknet_leaf_50_clk),
    .D(net34),
    .Q(net700));
 sky130_fd_sc_hd__dfxtp_1 s893 (.CLK(clknet_leaf_48_clk),
    .D(net43),
    .Q(net701));
 sky130_fd_sc_hd__dfxtp_1 s894 (.CLK(clknet_leaf_48_clk),
    .D(net44),
    .Q(net702));
 sky130_fd_sc_hd__dlclkp_1 s895 (.CLK(clknet_leaf_47_clk),
    .GATE(net56),
    .GCLK(net703));
 sky130_fd_sc_hd__dlclkp_2 s896 (.CLK(clknet_leaf_47_clk),
    .GATE(net57),
    .GCLK(net704));
 sky130_fd_sc_hd__dlclkp_4 s897 (.CLK(clknet_leaf_45_clk),
    .GATE(net61),
    .GCLK(net705));
 sky130_fd_sc_hd__dlxbn_2 s898 (.D(net62),
    .GATE_N(clknet_leaf_46_clk),
    .Q(net707),
    .Q_N(net706));
 sky130_fd_sc_hd__dlxbn_1 s899 (.D(net67),
    .GATE_N(clknet_leaf_2_clk),
    .Q(net709),
    .Q_N(net708));
 sky130_fd_sc_hd__dlxbp_1 s900 (.D(net68),
    .GATE(clknet_leaf_37_clk),
    .Q(net711),
    .Q_N(net710));
 sky130_fd_sc_hd__dlxtn_4 s901 (.D(net69),
    .GATE_N(clknet_leaf_44_clk),
    .Q(net712));
 sky130_fd_sc_hd__dlxtn_2 s902 (.D(net71),
    .GATE_N(clknet_leaf_44_clk),
    .Q(net713));
 sky130_fd_sc_hd__dlxtn_4 s903 (.D(net75),
    .GATE_N(clknet_leaf_44_clk),
    .Q(net714));
 sky130_fd_sc_hd__dlxtp_1 s904 (.D(net84),
    .GATE(clknet_leaf_45_clk),
    .Q(net715));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s905 (.D(net86),
    .SLEEP_B(clknet_leaf_39_clk),
    .Q(net716));
 sky130_fd_sc_hd__dfxbp_1 s906 (.CLK(clknet_leaf_39_clk),
    .D(net90),
    .Q(net718),
    .Q_N(net717));
 sky130_fd_sc_hd__dfxbp_2 s907 (.CLK(clknet_leaf_38_clk),
    .D(net91),
    .Q(net720),
    .Q_N(net719));
 sky130_fd_sc_hd__dfxtp_4 s908 (.CLK(clknet_leaf_38_clk),
    .D(net92),
    .Q(net721));
 sky130_fd_sc_hd__dfxtp_2 s909 (.CLK(clknet_leaf_41_clk),
    .D(net93),
    .Q(net722));
 sky130_fd_sc_hd__dfxtp_1 s910 (.CLK(clknet_leaf_38_clk),
    .D(net94),
    .Q(net723));
 sky130_fd_sc_hd__dlclkp_1 s911 (.CLK(clknet_leaf_39_clk),
    .GATE(net95),
    .GCLK(net724));
 sky130_fd_sc_hd__dlclkp_2 s912 (.CLK(clknet_leaf_38_clk),
    .GATE(net96),
    .GCLK(net725));
 sky130_fd_sc_hd__dlclkp_4 s913 (.CLK(clknet_leaf_37_clk),
    .GATE(net97),
    .GCLK(net726));
 sky130_fd_sc_hd__dlxbn_2 s914 (.D(net98),
    .GATE_N(clknet_leaf_39_clk),
    .Q(net728),
    .Q_N(net727));
 sky130_fd_sc_hd__dlxbn_1 s915 (.D(net99),
    .GATE_N(clknet_leaf_37_clk),
    .Q(net730),
    .Q_N(net729));
 sky130_fd_sc_hd__dlxbp_1 s916 (.D(net105),
    .GATE(clknet_leaf_41_clk),
    .Q(net1001),
    .Q_N(net731));
 sky130_fd_sc_hd__dlxtn_1 s917 (.D(net106),
    .GATE_N(clknet_leaf_38_clk),
    .Q(net732));
 sky130_fd_sc_hd__dlxtn_1 s918 (.D(net108),
    .GATE_N(clknet_leaf_38_clk),
    .Q(net733));
 sky130_fd_sc_hd__dlxtn_2 s919 (.D(net111),
    .GATE_N(clknet_leaf_37_clk),
    .Q(net734));
 sky130_fd_sc_hd__dlxtp_1 s920 (.D(net114),
    .GATE(clknet_leaf_37_clk),
    .Q(net735));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s921 (.D(net115),
    .SLEEP_B(clknet_leaf_33_clk),
    .Q(net736));
 sky130_fd_sc_hd__dfxbp_1 s922 (.CLK(clknet_leaf_37_clk),
    .D(net116),
    .Q(net738),
    .Q_N(net737));
 sky130_fd_sc_hd__dfxbp_1 s923 (.CLK(clknet_leaf_34_clk),
    .D(net118),
    .Q(net995),
    .Q_N(net739));
 sky130_fd_sc_hd__dfxtp_1 s924 (.CLK(clknet_leaf_34_clk),
    .D(net120),
    .Q(net740));
 sky130_fd_sc_hd__dfxtp_2 s925 (.CLK(clknet_leaf_34_clk),
    .D(net122),
    .Q(net741));
 sky130_fd_sc_hd__dfxtp_1 s926 (.CLK(clknet_leaf_36_clk),
    .D(net128),
    .Q(net742));
 sky130_fd_sc_hd__dlclkp_1 s927 (.CLK(clknet_leaf_1_clk),
    .GATE(net155),
    .GCLK(net743));
 sky130_fd_sc_hd__dlclkp_2 s928 (.CLK(clknet_leaf_1_clk),
    .GATE(net156),
    .GCLK(net744));
 sky130_fd_sc_hd__dlclkp_4 s929 (.CLK(clknet_leaf_1_clk),
    .GATE(net157),
    .GCLK(net745));
 sky130_fd_sc_hd__dlxbn_2 s930 (.D(net159),
    .GATE_N(clknet_leaf_1_clk),
    .Q(net747),
    .Q_N(net746));
 sky130_fd_sc_hd__dlxbn_2 s931 (.D(net170),
    .GATE_N(clknet_leaf_43_clk),
    .Q(net749),
    .Q_N(net748));
 sky130_fd_sc_hd__dlxbp_1 s932 (.D(net171),
    .GATE(clknet_leaf_43_clk),
    .Q(net751),
    .Q_N(net750));
 sky130_fd_sc_hd__dlxtn_4 s933 (.D(net173),
    .GATE_N(clknet_leaf_43_clk),
    .Q(net752));
 sky130_fd_sc_hd__dlxtn_2 s934 (.D(net174),
    .GATE_N(clknet_leaf_1_clk),
    .Q(net753));
 sky130_fd_sc_hd__dlxtn_2 s935 (.D(net177),
    .GATE_N(clknet_leaf_2_clk),
    .Q(net754));
 sky130_fd_sc_hd__dlxtp_1 s936 (.D(net178),
    .GATE(clknet_leaf_2_clk),
    .Q(net755));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s937 (.D(net184),
    .SLEEP_B(clknet_leaf_3_clk),
    .Q(net756));
 sky130_fd_sc_hd__dfxbp_1 s938 (.CLK(clknet_leaf_3_clk),
    .D(net186),
    .Q(net758),
    .Q_N(net757));
 sky130_fd_sc_hd__dfxbp_2 s939 (.CLK(clknet_leaf_44_clk),
    .D(net190),
    .Q(net760),
    .Q_N(net759));
 sky130_fd_sc_hd__dfxtp_2 s940 (.CLK(clknet_leaf_42_clk),
    .D(net192),
    .Q(net761));
 sky130_fd_sc_hd__dfxtp_4 s941 (.CLK(clknet_leaf_41_clk),
    .D(net198),
    .Q(net762));
 sky130_fd_sc_hd__dfxtp_2 s942 (.CLK(clknet_leaf_42_clk),
    .D(net199),
    .Q(net763));
 sky130_fd_sc_hd__dlclkp_1 s943 (.CLK(clknet_leaf_39_clk),
    .GATE(net200),
    .GCLK(net764));
 sky130_fd_sc_hd__dlclkp_2 s944 (.CLK(clknet_leaf_39_clk),
    .GATE(net201),
    .GCLK(net765));
 sky130_fd_sc_hd__dlclkp_4 s945 (.CLK(clknet_leaf_41_clk),
    .GATE(net208),
    .GCLK(net766));
 sky130_fd_sc_hd__dlxbn_1 s946 (.D(net212),
    .GATE_N(clknet_leaf_30_clk),
    .Q(net1013),
    .Q_N(net767));
 sky130_fd_sc_hd__dlxbn_1 s947 (.D(net218),
    .GATE_N(clknet_leaf_41_clk),
    .Q(net769),
    .Q_N(net768));
 sky130_fd_sc_hd__dlxbp_1 s948 (.D(net220),
    .GATE(clknet_leaf_30_clk),
    .Q(net771),
    .Q_N(net770));
 sky130_fd_sc_hd__dlxtn_2 s949 (.D(net221),
    .GATE_N(clknet_leaf_30_clk),
    .Q(net1007));
 sky130_fd_sc_hd__dlxtn_4 s950 (.D(net224),
    .GATE_N(clknet_leaf_40_clk),
    .Q(net772));
 sky130_fd_sc_hd__dlxtn_2 s951 (.D(net229),
    .GATE_N(clknet_leaf_32_clk),
    .Q(net773));
 sky130_fd_sc_hd__dlxtp_1 s952 (.D(net231),
    .GATE(clknet_leaf_33_clk),
    .Q(net1005));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s953 (.D(net240),
    .SLEEP_B(clknet_leaf_30_clk),
    .Q(net774));
 sky130_fd_sc_hd__dfxbp_1 s954 (.CLK(clknet_leaf_31_clk),
    .D(net242),
    .Q(net776),
    .Q_N(net775));
 sky130_fd_sc_hd__dfxbp_1 s955 (.CLK(clknet_leaf_32_clk),
    .D(net245),
    .Q(net778),
    .Q_N(net777));
 sky130_fd_sc_hd__dfxtp_1 s956 (.CLK(clknet_leaf_8_clk),
    .D(net270),
    .Q(net779));
 sky130_fd_sc_hd__dfxtp_4 s957 (.CLK(clknet_leaf_8_clk),
    .D(net271),
    .Q(net780));
 sky130_fd_sc_hd__dfxtp_1 s958 (.CLK(clknet_leaf_7_clk),
    .D(net272),
    .Q(net781));
 sky130_fd_sc_hd__dlclkp_1 s959 (.CLK(clknet_leaf_3_clk),
    .GATE(net278),
    .GCLK(net782));
 sky130_fd_sc_hd__dlclkp_2 s960 (.CLK(clknet_leaf_5_clk),
    .GATE(net280),
    .GCLK(net783));
 sky130_fd_sc_hd__dlclkp_4 s961 (.CLK(clknet_leaf_3_clk),
    .GATE(net286),
    .GCLK(net784));
 sky130_fd_sc_hd__dlxbn_2 s962 (.D(net294),
    .GATE_N(clknet_leaf_5_clk),
    .Q(net786),
    .Q_N(net785));
 sky130_fd_sc_hd__dlxbn_2 s963 (.D(net297),
    .GATE_N(clknet_leaf_4_clk),
    .Q(net978),
    .Q_N(net787));
 sky130_fd_sc_hd__dlxbp_1 s964 (.D(net299),
    .GATE(clknet_leaf_4_clk),
    .Q(net789),
    .Q_N(net788));
 sky130_fd_sc_hd__dlxtn_2 s965 (.D(net304),
    .GATE_N(clknet_leaf_41_clk),
    .Q(net790));
 sky130_fd_sc_hd__dlxtn_1 s966 (.D(net305),
    .GATE_N(clknet_leaf_1_clk),
    .Q(net791));
 sky130_fd_sc_hd__dlxtn_2 s967 (.D(net307),
    .GATE_N(clknet_leaf_42_clk),
    .Q(net792));
 sky130_fd_sc_hd__dlxtp_1 s968 (.D(net308),
    .GATE(clknet_leaf_41_clk),
    .Q(net793));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s969 (.D(net310),
    .SLEEP_B(clknet_leaf_18_clk),
    .Q(net1011));
 sky130_fd_sc_hd__dfxbp_1 s970 (.CLK(clknet_leaf_29_clk),
    .D(net311),
    .Q(net795),
    .Q_N(net794));
 sky130_fd_sc_hd__dfxbp_2 s971 (.CLK(clknet_leaf_29_clk),
    .D(net314),
    .Q(net797),
    .Q_N(net796));
 sky130_fd_sc_hd__dfxtp_1 s972 (.CLK(clknet_leaf_29_clk),
    .D(net316),
    .Q(net798));
 sky130_fd_sc_hd__dfxtp_2 s973 (.CLK(clknet_leaf_18_clk),
    .D(net317),
    .Q(net1015));
 sky130_fd_sc_hd__dfxtp_1 s974 (.CLK(clknet_leaf_18_clk),
    .D(net318),
    .Q(net799));
 sky130_fd_sc_hd__dlclkp_1 s975 (.CLK(clknet_leaf_29_clk),
    .GATE(net319),
    .GCLK(net800));
 sky130_fd_sc_hd__dlclkp_2 s976 (.CLK(clknet_leaf_28_clk),
    .GATE(net323),
    .GCLK(net801));
 sky130_fd_sc_hd__dlclkp_4 s977 (.CLK(clknet_leaf_27_clk),
    .GATE(net329),
    .GCLK(net802));
 sky130_fd_sc_hd__dlxbn_1 s978 (.D(net330),
    .GATE_N(clknet_leaf_28_clk),
    .Q(net804),
    .Q_N(net803));
 sky130_fd_sc_hd__dlxbn_1 s979 (.D(net335),
    .GATE_N(clknet_leaf_28_clk),
    .Q(net975),
    .Q_N(net805));
 sky130_fd_sc_hd__dlxbp_1 s980 (.D(net337),
    .GATE(clknet_leaf_26_clk),
    .Q(net985),
    .Q_N(net806));
 sky130_fd_sc_hd__dlxtn_1 s981 (.D(net339),
    .GATE_N(clknet_leaf_26_clk),
    .Q(net807));
 sky130_fd_sc_hd__dlxtn_2 s982 (.D(net343),
    .GATE_N(clknet_leaf_30_clk),
    .Q(net808));
 sky130_fd_sc_hd__dlxtn_1 s983 (.D(net357),
    .GATE_N(clknet_leaf_32_clk),
    .Q(net809));
 sky130_fd_sc_hd__dlxtp_1 s984 (.D(net360),
    .GATE(clknet_leaf_25_clk),
    .Q(net810));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s985 (.D(net362),
    .SLEEP_B(clknet_leaf_24_clk),
    .Q(net811));
 sky130_fd_sc_hd__dfxbp_1 s986 (.CLK(clknet_leaf_32_clk),
    .D(net363),
    .Q(net1010),
    .Q_N(net812));
 sky130_fd_sc_hd__dfxbp_1 s987 (.CLK(clknet_leaf_10_clk),
    .D(net372),
    .Q(net814),
    .Q_N(net813));
 sky130_fd_sc_hd__dfxtp_1 s988 (.CLK(clknet_leaf_9_clk),
    .D(net379),
    .Q(net815));
 sky130_fd_sc_hd__dfxtp_2 s989 (.CLK(clknet_leaf_10_clk),
    .D(net383),
    .Q(net816));
 sky130_fd_sc_hd__dfxtp_2 s990 (.CLK(clknet_leaf_9_clk),
    .D(net384),
    .Q(net817));
 sky130_fd_sc_hd__dlclkp_1 s991 (.CLK(clknet_leaf_10_clk),
    .GATE(net386),
    .GCLK(net818));
 sky130_fd_sc_hd__dlclkp_2 s992 (.CLK(clknet_leaf_10_clk),
    .GATE(net388),
    .GCLK(net819));
 sky130_fd_sc_hd__dlclkp_4 s993 (.CLK(clknet_leaf_9_clk),
    .GATE(net392),
    .GCLK(net820));
 sky130_fd_sc_hd__dlxbn_1 s994 (.D(net401),
    .GATE_N(clknet_leaf_16_clk),
    .Q(net822),
    .Q_N(net821));
 sky130_fd_sc_hd__dlxbn_1 s995 (.D(net403),
    .GATE_N(clknet_leaf_10_clk),
    .Q(net824),
    .Q_N(net823));
 sky130_fd_sc_hd__dlxbp_1 s996 (.D(net405),
    .GATE(clknet_leaf_16_clk),
    .Q(net826),
    .Q_N(net825));
 sky130_fd_sc_hd__dlxtn_2 s997 (.D(net408),
    .GATE_N(clknet_leaf_15_clk),
    .Q(net827));
 sky130_fd_sc_hd__dlxtn_1 s998 (.D(net409),
    .GATE_N(clknet_leaf_15_clk),
    .Q(net828));
 sky130_fd_sc_hd__dlxtn_2 s999 (.D(net411),
    .GATE_N(clknet_leaf_16_clk),
    .Q(net829));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(in0),
    .X(net412));
 sky130_fd_sc_hd__buf_1 input2 (.A(in1),
    .X(net869));
 sky130_fd_sc_hd__buf_2 input3 (.A(in10),
    .X(net870));
 sky130_fd_sc_hd__buf_2 input4 (.A(in11),
    .X(net871));
 sky130_fd_sc_hd__buf_1 input5 (.A(in12),
    .X(net872));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(in13),
    .X(net873));
 sky130_fd_sc_hd__buf_2 input7 (.A(in14),
    .X(net874));
 sky130_fd_sc_hd__buf_2 input8 (.A(in15),
    .X(net875));
 sky130_fd_sc_hd__buf_1 input9 (.A(in16),
    .X(net876));
 sky130_fd_sc_hd__buf_2 input10 (.A(in17),
    .X(net877));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(in18),
    .X(net878));
 sky130_fd_sc_hd__buf_1 input12 (.A(in19),
    .X(net879));
 sky130_fd_sc_hd__buf_2 input13 (.A(in2),
    .X(net880));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(in20),
    .X(net881));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(in21),
    .X(net882));
 sky130_fd_sc_hd__buf_2 input16 (.A(in22),
    .X(net883));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(in23),
    .X(net884));
 sky130_fd_sc_hd__buf_1 input18 (.A(in24),
    .X(net885));
 sky130_fd_sc_hd__buf_1 input19 (.A(in25),
    .X(net886));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(in26),
    .X(net887));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(in27),
    .X(net888));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(in28),
    .X(net889));
 sky130_fd_sc_hd__clkbuf_4 input23 (.A(in29),
    .X(net890));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(in3),
    .X(net891));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(in30),
    .X(net892));
 sky130_fd_sc_hd__clkbuf_4 input26 (.A(in31),
    .X(net893));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(in32),
    .X(net894));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(in33),
    .X(net895));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(in34),
    .X(net896));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(in35),
    .X(net897));
 sky130_fd_sc_hd__buf_2 input31 (.A(in36),
    .X(net898));
 sky130_fd_sc_hd__buf_1 input32 (.A(in37),
    .X(net899));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(in38),
    .X(net900));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(in39),
    .X(net901));
 sky130_fd_sc_hd__buf_2 input35 (.A(in4),
    .X(net902));
 sky130_fd_sc_hd__clkbuf_8 input36 (.A(in40),
    .X(net903));
 sky130_fd_sc_hd__buf_4 input37 (.A(in41),
    .X(net904));
 sky130_fd_sc_hd__buf_2 input38 (.A(in42),
    .X(net905));
 sky130_fd_sc_hd__buf_4 input39 (.A(in43),
    .X(net906));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(in44),
    .X(net907));
 sky130_fd_sc_hd__clkbuf_4 input41 (.A(in45),
    .X(net908));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(in46),
    .X(net909));
 sky130_fd_sc_hd__buf_1 input43 (.A(in47),
    .X(net910));
 sky130_fd_sc_hd__clkbuf_4 input44 (.A(in48),
    .X(net911));
 sky130_fd_sc_hd__buf_1 input45 (.A(in49),
    .X(net912));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(in5),
    .X(net913));
 sky130_fd_sc_hd__buf_1 input47 (.A(in50),
    .X(net914));
 sky130_fd_sc_hd__buf_2 input48 (.A(in51),
    .X(net915));
 sky130_fd_sc_hd__clkbuf_4 input49 (.A(in52),
    .X(net916));
 sky130_fd_sc_hd__clkbuf_4 input50 (.A(in53),
    .X(net917));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(in54),
    .X(net918));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(in55),
    .X(net919));
 sky130_fd_sc_hd__clkbuf_8 input53 (.A(in56),
    .X(net920));
 sky130_fd_sc_hd__buf_2 input54 (.A(in57),
    .X(net921));
 sky130_fd_sc_hd__buf_4 input55 (.A(in58),
    .X(net922));
 sky130_fd_sc_hd__buf_1 input56 (.A(in59),
    .X(net923));
 sky130_fd_sc_hd__dlymetal6s2s_1 input57 (.A(in6),
    .X(net924));
 sky130_fd_sc_hd__buf_2 input58 (.A(in60),
    .X(net925));
 sky130_fd_sc_hd__buf_2 input59 (.A(in61),
    .X(net926));
 sky130_fd_sc_hd__buf_4 input60 (.A(in62),
    .X(net927));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(in63),
    .X(net928));
 sky130_fd_sc_hd__buf_2 input62 (.A(in64),
    .X(net929));
 sky130_fd_sc_hd__dlymetal6s2s_1 input63 (.A(in65),
    .X(net930));
 sky130_fd_sc_hd__buf_1 input64 (.A(in66),
    .X(net931));
 sky130_fd_sc_hd__buf_1 input65 (.A(in67),
    .X(net932));
 sky130_fd_sc_hd__buf_1 input66 (.A(in68),
    .X(net933));
 sky130_fd_sc_hd__clkbuf_4 input67 (.A(in69),
    .X(net934));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(in7),
    .X(net935));
 sky130_fd_sc_hd__clkbuf_4 input69 (.A(in70),
    .X(net936));
 sky130_fd_sc_hd__buf_1 input70 (.A(in71),
    .X(net937));
 sky130_fd_sc_hd__buf_2 input71 (.A(in72),
    .X(net938));
 sky130_fd_sc_hd__clkbuf_2 input72 (.A(in73),
    .X(net939));
 sky130_fd_sc_hd__clkbuf_4 input73 (.A(in74),
    .X(net940));
 sky130_fd_sc_hd__clkbuf_4 input74 (.A(in75),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_2 input75 (.A(in76),
    .X(net942));
 sky130_fd_sc_hd__buf_1 input76 (.A(in77),
    .X(net943));
 sky130_fd_sc_hd__buf_1 input77 (.A(in78),
    .X(net944));
 sky130_fd_sc_hd__buf_1 input78 (.A(in79),
    .X(net945));
 sky130_fd_sc_hd__buf_1 input79 (.A(in8),
    .X(net946));
 sky130_fd_sc_hd__buf_1 input80 (.A(in80),
    .X(net947));
 sky130_fd_sc_hd__buf_1 input81 (.A(in81),
    .X(net948));
 sky130_fd_sc_hd__clkbuf_4 input82 (.A(in82),
    .X(net949));
 sky130_fd_sc_hd__buf_2 input83 (.A(in83),
    .X(net950));
 sky130_fd_sc_hd__buf_1 input84 (.A(in84),
    .X(net951));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(in85),
    .X(net952));
 sky130_fd_sc_hd__buf_1 input86 (.A(in86),
    .X(net953));
 sky130_fd_sc_hd__buf_1 input87 (.A(in87),
    .X(net954));
 sky130_fd_sc_hd__buf_1 input88 (.A(in88),
    .X(net955));
 sky130_fd_sc_hd__buf_1 input89 (.A(in89),
    .X(net956));
 sky130_fd_sc_hd__clkbuf_2 input90 (.A(in9),
    .X(net957));
 sky130_fd_sc_hd__buf_1 input91 (.A(in90),
    .X(net958));
 sky130_fd_sc_hd__clkbuf_4 input92 (.A(in91),
    .X(net959));
 sky130_fd_sc_hd__clkbuf_4 input93 (.A(in92),
    .X(net960));
 sky130_fd_sc_hd__buf_4 input94 (.A(in93),
    .X(net961));
 sky130_fd_sc_hd__buf_2 input95 (.A(in94),
    .X(net962));
 sky130_fd_sc_hd__buf_1 input96 (.A(in95),
    .X(net963));
 sky130_fd_sc_hd__buf_1 input97 (.A(in96),
    .X(net964));
 sky130_fd_sc_hd__buf_2 input98 (.A(in97),
    .X(net965));
 sky130_fd_sc_hd__dlymetal6s2s_1 input99 (.A(in98),
    .X(net966));
 sky130_fd_sc_hd__buf_1 input100 (.A(in99),
    .X(net967));
 sky130_fd_sc_hd__buf_2 output101 (.A(net1060),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(clknet_1_1__leaf_net969),
    .X(out10));
 sky130_fd_sc_hd__clkbuf_1 output103 (.A(clknet_1_1__leaf_net970),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net971),
    .X(out12));
 sky130_fd_sc_hd__clkbuf_4 output105 (.A(net1063),
    .X(out13));
 sky130_fd_sc_hd__clkbuf_4 output106 (.A(net973),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output107 (.A(net974),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output108 (.A(net975),
    .X(out18));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(clknet_1_1__leaf_net976),
    .X(out19));
 sky130_fd_sc_hd__clkbuf_4 output110 (.A(net977),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output111 (.A(net978),
    .X(out20));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(clknet_1_1__leaf_net979),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_4 output113 (.A(net980),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output114 (.A(net981),
    .X(out24));
 sky130_fd_sc_hd__clkbuf_4 output115 (.A(net982),
    .X(out25));
 sky130_fd_sc_hd__buf_2 output116 (.A(net983),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output117 (.A(net984),
    .X(out27));
 sky130_fd_sc_hd__buf_2 output118 (.A(net985),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output119 (.A(net986),
    .X(out29));
 sky130_fd_sc_hd__clkbuf_1 output120 (.A(clknet_1_1__leaf_net987),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output121 (.A(net988),
    .X(out31));
 sky130_fd_sc_hd__clkbuf_4 output122 (.A(net989),
    .X(out32));
 sky130_fd_sc_hd__clkbuf_1 output123 (.A(clknet_1_1__leaf_net990),
    .X(out33));
 sky130_fd_sc_hd__buf_2 output124 (.A(net991),
    .X(out34));
 sky130_fd_sc_hd__clkbuf_1 output125 (.A(clknet_1_1__leaf_net992),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output126 (.A(net993),
    .X(out36));
 sky130_fd_sc_hd__buf_2 output127 (.A(net994),
    .X(out37));
 sky130_fd_sc_hd__buf_2 output128 (.A(net995),
    .X(out38));
 sky130_fd_sc_hd__clkbuf_1 output129 (.A(clknet_1_1__leaf_net996),
    .X(out39));
 sky130_fd_sc_hd__buf_2 output130 (.A(net997),
    .X(out42));
 sky130_fd_sc_hd__clkbuf_1 output131 (.A(net998),
    .X(out43));
 sky130_fd_sc_hd__clkbuf_1 output132 (.A(clknet_1_1__leaf_net999),
    .X(out45));
 sky130_fd_sc_hd__clkbuf_1 output133 (.A(clknet_1_1__leaf_net1000),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output134 (.A(net1001),
    .X(out48));
 sky130_fd_sc_hd__clkbuf_1 output135 (.A(clknet_1_0__leaf_net1002),
    .X(out49));
 sky130_fd_sc_hd__clkbuf_1 output136 (.A(clknet_1_1__leaf_net1003),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output137 (.A(net1004),
    .X(out51));
 sky130_fd_sc_hd__buf_2 output138 (.A(net1005),
    .X(out52));
 sky130_fd_sc_hd__buf_2 output139 (.A(net1006),
    .X(out53));
 sky130_fd_sc_hd__buf_2 output140 (.A(net1007),
    .X(out54));
 sky130_fd_sc_hd__buf_2 output141 (.A(net1008),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output142 (.A(net1009),
    .X(out57));
 sky130_fd_sc_hd__buf_2 output143 (.A(net1010),
    .X(out58));
 sky130_fd_sc_hd__buf_2 output144 (.A(net1011),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output145 (.A(net1012),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output146 (.A(net1013),
    .X(out60));
 sky130_fd_sc_hd__buf_2 output147 (.A(net1014),
    .X(out62));
 sky130_fd_sc_hd__buf_2 output148 (.A(net1015),
    .X(out63));
 sky130_fd_sc_hd__buf_2 output149 (.A(net1016),
    .X(out64));
 sky130_fd_sc_hd__buf_2 output150 (.A(net1017),
    .X(out66));
 sky130_fd_sc_hd__buf_2 output151 (.A(net1018),
    .X(out67));
 sky130_fd_sc_hd__buf_2 output152 (.A(net1019),
    .X(out68));
 sky130_fd_sc_hd__buf_2 output153 (.A(net1020),
    .X(out69));
 sky130_fd_sc_hd__buf_2 output154 (.A(net1021),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_1 output155 (.A(clknet_1_1__leaf_net1022),
    .X(out70));
 sky130_fd_sc_hd__buf_2 output156 (.A(net1023),
    .X(out71));
 sky130_fd_sc_hd__buf_2 output157 (.A(net1024),
    .X(out73));
 sky130_fd_sc_hd__buf_2 output158 (.A(net1025),
    .X(out75));
 sky130_fd_sc_hd__buf_2 output159 (.A(net1026),
    .X(out76));
 sky130_fd_sc_hd__buf_2 output160 (.A(net1027),
    .X(out77));
 sky130_fd_sc_hd__buf_2 output161 (.A(net1028),
    .X(out78));
 sky130_fd_sc_hd__buf_2 output162 (.A(net1029),
    .X(out79));
 sky130_fd_sc_hd__clkbuf_1 output163 (.A(net1030),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output164 (.A(net1031),
    .X(out80));
 sky130_fd_sc_hd__buf_2 output165 (.A(net1032),
    .X(out81));
 sky130_fd_sc_hd__buf_2 output166 (.A(net1033),
    .X(out82));
 sky130_fd_sc_hd__buf_2 output167 (.A(net1034),
    .X(out84));
 sky130_fd_sc_hd__buf_2 output168 (.A(net1035),
    .X(out85));
 sky130_fd_sc_hd__buf_2 output169 (.A(net1036),
    .X(out86));
 sky130_fd_sc_hd__buf_2 output170 (.A(net1037),
    .X(out87));
 sky130_fd_sc_hd__buf_2 output171 (.A(net1038),
    .X(out88));
 sky130_fd_sc_hd__buf_2 output172 (.A(net1039),
    .X(out89));
 sky130_fd_sc_hd__buf_2 output173 (.A(net1040),
    .X(out9));
 sky130_fd_sc_hd__buf_2 output174 (.A(net1041),
    .X(out90));
 sky130_fd_sc_hd__buf_2 output175 (.A(net1042),
    .X(out91));
 sky130_fd_sc_hd__buf_2 output176 (.A(net1043),
    .X(out93));
 sky130_fd_sc_hd__buf_2 output177 (.A(net1044),
    .X(out94));
 sky130_fd_sc_hd__buf_2 output178 (.A(net1045),
    .X(out95));
 sky130_fd_sc_hd__buf_2 output179 (.A(net1046),
    .X(out96));
 sky130_fd_sc_hd__buf_2 output180 (.A(net1047),
    .X(out97));
 sky130_fd_sc_hd__buf_2 output181 (.A(net1048),
    .X(out99));
 sky130_fd_sc_hd__clkbuf_4 fanout182 (.A(net247),
    .X(net1049));
 sky130_fd_sc_hd__buf_2 fanout183 (.A(net1052),
    .X(net1050));
 sky130_fd_sc_hd__clkbuf_4 fanout184 (.A(net1052),
    .X(net1051));
 sky130_fd_sc_hd__clkbuf_4 fanout185 (.A(net154),
    .X(net1052));
 sky130_fd_sc_hd__buf_4 fanout186 (.A(net146),
    .X(net1053));
 sky130_fd_sc_hd__clkbuf_4 fanout187 (.A(net55),
    .X(net1054));
 sky130_fd_sc_hd__buf_4 fanout188 (.A(net53),
    .X(net1055));
 sky130_fd_sc_hd__buf_4 fanout189 (.A(net41),
    .X(net1056));
 sky130_fd_sc_hd__buf_4 fanout190 (.A(net37),
    .X(net1057));
 sky130_fd_sc_hd__buf_4 fanout191 (.A(net27),
    .X(net1058));
 sky130_fd_sc_hd__clkbuf_2 fanout192 (.A(net27),
    .X(net1059));
 sky130_fd_sc_hd__buf_4 fanout193 (.A(net968),
    .X(net1060));
 sky130_fd_sc_hd__clkbuf_4 fanout194 (.A(net968),
    .X(net1061));
 sky130_fd_sc_hd__buf_2 fanout195 (.A(net1063),
    .X(net1062));
 sky130_fd_sc_hd__clkbuf_4 fanout196 (.A(net972),
    .X(net1063));
 sky130_fd_sc_hd__clkbuf_4 fanout197 (.A(net195),
    .X(net1064));
 sky130_fd_sc_hd__clkbuf_2 fanout198 (.A(net195),
    .X(net1065));
 sky130_fd_sc_hd__buf_2 fanout199 (.A(net1067),
    .X(net1066));
 sky130_fd_sc_hd__clkbuf_2 fanout200 (.A(net1068),
    .X(net1067));
 sky130_fd_sc_hd__clkbuf_2 fanout201 (.A(net1069),
    .X(net1068));
 sky130_fd_sc_hd__clkbuf_4 fanout202 (.A(net134),
    .X(net1069));
 sky130_fd_sc_hd__buf_4 fanout203 (.A(net65),
    .X(net1070));
 sky130_fd_sc_hd__clkbuf_4 fanout204 (.A(net1072),
    .X(net1071));
 sky130_fd_sc_hd__clkbuf_4 fanout205 (.A(net50),
    .X(net1072));
 sky130_fd_sc_hd__buf_4 fanout206 (.A(net26),
    .X(net1073));
 sky130_fd_sc_hd__clkbuf_4 fanout207 (.A(net23),
    .X(net1074));
 sky130_fd_sc_hd__clkbuf_4 fanout208 (.A(net774),
    .X(net1075));
 sky130_fd_sc_hd__clkbuf_4 wire209 (.A(net755),
    .X(net1076));
 sky130_fd_sc_hd__buf_4 fanout210 (.A(net733),
    .X(net1077));
 sky130_fd_sc_hd__buf_4 max_cap211 (.A(net716),
    .X(net1078));
 sky130_fd_sc_hd__buf_2 max_cap212 (.A(net715),
    .X(net1079));
 sky130_fd_sc_hd__buf_4 fanout213 (.A(net702),
    .X(net1080));
 sky130_fd_sc_hd__clkbuf_2 fanout214 (.A(net702),
    .X(net1081));
 sky130_fd_sc_hd__clkbuf_8 fanout215 (.A(net701),
    .X(net1082));
 sky130_fd_sc_hd__buf_2 fanout216 (.A(net701),
    .X(net1083));
 sky130_fd_sc_hd__clkbuf_4 max_cap217 (.A(net831),
    .X(net1084));
 sky130_fd_sc_hd__buf_2 max_cap218 (.A(net598),
    .X(net1085));
 sky130_fd_sc_hd__clkbuf_4 fanout219 (.A(net142),
    .X(net1086));
 sky130_fd_sc_hd__buf_4 fanout220 (.A(net143),
    .X(net1087));
 sky130_fd_sc_hd__clkbuf_2 max_cap221 (.A(net42),
    .X(net1088));
 sky130_fd_sc_hd__buf_4 max_cap222 (.A(net983),
    .X(net1089));
 sky130_fd_sc_hd__clkbuf_4 fanout223 (.A(net28),
    .X(net1090));
 sky130_fd_sc_hd__clkbuf_4 fanout224 (.A(net29),
    .X(net1091));
 sky130_fd_sc_hd__buf_4 fanout225 (.A(net1039),
    .X(net1092));
 sky130_fd_sc_hd__buf_4 fanout226 (.A(net957),
    .X(net1093));
 sky130_fd_sc_hd__clkbuf_4 fanout227 (.A(net876),
    .X(net1094));
 sky130_fd_sc_hd__buf_4 fanout228 (.A(net875),
    .X(net1095));
 sky130_fd_sc_hd__clkbuf_2 fanout229 (.A(net875),
    .X(net1096));
 sky130_fd_sc_hd__buf_4 fanout230 (.A(net1098),
    .X(net1097));
 sky130_fd_sc_hd__buf_4 fanout231 (.A(net946),
    .X(net1098));
 sky130_fd_sc_hd__clkbuf_8 fanout232 (.A(net874),
    .X(net1099));
 sky130_fd_sc_hd__buf_4 fanout233 (.A(net935),
    .X(net1100));
 sky130_fd_sc_hd__clkbuf_2 fanout234 (.A(net935),
    .X(net1101));
 sky130_fd_sc_hd__buf_4 fanout235 (.A(net924),
    .X(net1102));
 sky130_fd_sc_hd__clkbuf_2 fanout236 (.A(net924),
    .X(net1103));
 sky130_fd_sc_hd__buf_4 fanout237 (.A(net872),
    .X(net1104));
 sky130_fd_sc_hd__buf_2 fanout238 (.A(net872),
    .X(net1105));
 sky130_fd_sc_hd__buf_4 fanout239 (.A(net913),
    .X(net1106));
 sky130_fd_sc_hd__buf_4 fanout240 (.A(net871),
    .X(net1107));
 sky130_fd_sc_hd__buf_4 fanout241 (.A(net902),
    .X(net1108));
 sky130_fd_sc_hd__buf_4 fanout242 (.A(net899),
    .X(net1109));
 sky130_fd_sc_hd__buf_4 fanout243 (.A(net892),
    .X(net1110));
 sky130_fd_sc_hd__clkbuf_4 fanout244 (.A(net1112),
    .X(net1111));
 sky130_fd_sc_hd__buf_2 fanout245 (.A(net1114),
    .X(net1112));
 sky130_fd_sc_hd__clkbuf_4 fanout246 (.A(net1114),
    .X(net1113));
 sky130_fd_sc_hd__buf_2 fanout247 (.A(net891),
    .X(net1114));
 sky130_fd_sc_hd__clkbuf_4 fanout248 (.A(net1116),
    .X(net1115));
 sky130_fd_sc_hd__clkbuf_4 fanout249 (.A(net891),
    .X(net1116));
 sky130_fd_sc_hd__buf_4 fanout250 (.A(net869),
    .X(net1117));
 sky130_fd_sc_hd__buf_4 fanout251 (.A(net886),
    .X(net1118));
 sky130_fd_sc_hd__buf_2 fanout252 (.A(net886),
    .X(net1119));
 sky130_fd_sc_hd__clkbuf_4 fanout253 (.A(net885),
    .X(net1120));
 sky130_fd_sc_hd__buf_4 fanout254 (.A(net882),
    .X(net1121));
 sky130_fd_sc_hd__buf_4 fanout255 (.A(net881),
    .X(net1122));
 sky130_fd_sc_hd__clkbuf_4 fanout256 (.A(net880),
    .X(net1123));
 sky130_fd_sc_hd__clkbuf_4 fanout257 (.A(net879),
    .X(net1124));
 sky130_fd_sc_hd__clkbuf_4 fanout258 (.A(net878),
    .X(net1125));
 sky130_fd_sc_hd__clkbuf_8 fanout259 (.A(net877),
    .X(net1126));
 sky130_fd_sc_hd__buf_4 fanout260 (.A(net412),
    .X(net1127));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_36_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_37_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_38_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_39_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_40_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_41_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_42_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_43_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_44_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_45_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_46_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_47_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_48_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_49_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_50_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net820 (.A(net820),
    .X(clknet_0_net820));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net820 (.A(clknet_0_net820),
    .X(clknet_1_0__leaf_net820));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net820 (.A(clknet_0_net820),
    .X(clknet_1_1__leaf_net820));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net529 (.A(net529),
    .X(clknet_0_net529));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net529 (.A(clknet_0_net529),
    .X(clknet_1_0__leaf_net529));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net529 (.A(clknet_0_net529),
    .X(clknet_1_1__leaf_net529));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net859 (.A(net859),
    .X(clknet_0_net859));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net859 (.A(clknet_0_net859),
    .X(clknet_1_0__leaf_net859));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net859 (.A(clknet_0_net859),
    .X(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net523 (.A(net523),
    .X(clknet_0_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net523 (.A(clknet_0_net523),
    .X(clknet_1_0__leaf_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net523 (.A(clknet_0_net523),
    .X(clknet_1_1__leaf_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net860 (.A(net860),
    .X(clknet_0_net860));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net860 (.A(clknet_0_net860),
    .X(clknet_1_0__leaf_net860));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net860 (.A(clknet_0_net860),
    .X(clknet_1_1__leaf_net860));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net539 (.A(net539),
    .X(clknet_0_net539));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net539 (.A(clknet_0_net539),
    .X(clknet_1_0__leaf_net539));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net539 (.A(clknet_0_net539),
    .X(clknet_1_1__leaf_net539));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net564 (.A(net564),
    .X(clknet_0_net564));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net564 (.A(clknet_0_net564),
    .X(clknet_1_0__leaf_net564));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net564 (.A(clknet_0_net564),
    .X(clknet_1_1__leaf_net564));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net681 (.A(net681),
    .X(clknet_0_net681));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net681 (.A(clknet_0_net681),
    .X(clknet_1_0__leaf_net681));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net681 (.A(clknet_0_net681),
    .X(clknet_1_1__leaf_net681));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net516 (.A(net516),
    .X(clknet_0_net516));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net516 (.A(clknet_0_net516),
    .X(clknet_1_0__leaf_net516));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net516 (.A(clknet_0_net516),
    .X(clknet_1_1__leaf_net516));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net992 (.A(net992),
    .X(clknet_0_net992));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net992 (.A(clknet_0_net992),
    .X(clknet_1_0__leaf_net992));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net992 (.A(clknet_0_net992),
    .X(clknet_1_1__leaf_net992));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net406 (.A(net406),
    .X(clknet_0_net406));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net406 (.A(clknet_0_net406),
    .X(clknet_1_0__leaf_net406));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net406 (.A(clknet_0_net406),
    .X(clknet_1_1__leaf_net406));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net651 (.A(net651),
    .X(clknet_0_net651));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net651 (.A(clknet_0_net651),
    .X(clknet_1_0__leaf_net651));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net651 (.A(clknet_0_net651),
    .X(clknet_1_1__leaf_net651));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net819 (.A(net819),
    .X(clknet_0_net819));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net819 (.A(clknet_0_net819),
    .X(clknet_1_0__leaf_net819));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net819 (.A(clknet_0_net819),
    .X(clknet_1_1__leaf_net819));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net391 (.A(net391),
    .X(clknet_0_net391));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net391 (.A(clknet_0_net391),
    .X(clknet_1_0__leaf_net391));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net391 (.A(clknet_0_net391),
    .X(clknet_1_1__leaf_net391));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net858 (.A(net858),
    .X(clknet_0_net858));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net858 (.A(clknet_0_net858),
    .X(clknet_1_0__leaf_net858));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net858 (.A(clknet_0_net858),
    .X(clknet_1_1__leaf_net858));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net818 (.A(net818),
    .X(clknet_0_net818));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net818 (.A(clknet_0_net818),
    .X(clknet_1_0__leaf_net818));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net818 (.A(clknet_0_net818),
    .X(clknet_1_1__leaf_net818));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net488 (.A(net488),
    .X(clknet_0_net488));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net488 (.A(clknet_0_net488),
    .X(clknet_1_0__leaf_net488));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net488 (.A(clknet_0_net488),
    .X(clknet_1_1__leaf_net488));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net394 (.A(net394),
    .X(clknet_0_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net394 (.A(clknet_0_net394),
    .X(clknet_1_0__leaf_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net394 (.A(clknet_0_net394),
    .X(clknet_1_1__leaf_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net393 (.A(net393),
    .X(clknet_0_net393));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net393 (.A(clknet_0_net393),
    .X(clknet_1_0__leaf_net393));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net393 (.A(clknet_0_net393),
    .X(clknet_1_1__leaf_net393));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net839 (.A(net839),
    .X(clknet_0_net839));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net839 (.A(clknet_0_net839),
    .X(clknet_1_0__leaf_net839));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net839 (.A(clknet_0_net839),
    .X(clknet_1_1__leaf_net839));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net464 (.A(net464),
    .X(clknet_0_net464));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net464 (.A(clknet_0_net464),
    .X(clknet_1_0__leaf_net464));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net464 (.A(clknet_0_net464),
    .X(clknet_1_1__leaf_net464));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net462 (.A(net462),
    .X(clknet_0_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net462 (.A(clknet_0_net462),
    .X(clknet_1_0__leaf_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net462 (.A(clknet_0_net462),
    .X(clknet_1_1__leaf_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net970 (.A(net970),
    .X(clknet_0_net970));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net970 (.A(clknet_0_net970),
    .X(clknet_1_0__leaf_net970));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net970 (.A(clknet_0_net970),
    .X(clknet_1_1__leaf_net970));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net390 (.A(net390),
    .X(clknet_0_net390));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net390 (.A(clknet_0_net390),
    .X(clknet_1_0__leaf_net390));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net390 (.A(clknet_0_net390),
    .X(clknet_1_1__leaf_net390));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net389 (.A(net389),
    .X(clknet_0_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_0__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_1__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net387 (.A(net387),
    .X(clknet_0_net387));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net387 (.A(clknet_0_net387),
    .X(clknet_1_0__leaf_net387));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net387 (.A(clknet_0_net387),
    .X(clknet_1_1__leaf_net387));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net802 (.A(net802),
    .X(clknet_0_net802));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net802 (.A(clknet_0_net802),
    .X(clknet_1_0__leaf_net802));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net802 (.A(clknet_0_net802),
    .X(clknet_1_1__leaf_net802));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1000 (.A(net1000),
    .X(clknet_0_net1000));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1000 (.A(clknet_0_net1000),
    .X(clknet_1_0__leaf_net1000));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1000 (.A(clknet_0_net1000),
    .X(clknet_1_1__leaf_net1000));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net341 (.A(net341),
    .X(clknet_0_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net341 (.A(clknet_0_net341),
    .X(clknet_1_0__leaf_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net341 (.A(clknet_0_net341),
    .X(clknet_1_1__leaf_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net332 (.A(net332),
    .X(clknet_0_net332));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net332 (.A(clknet_0_net332),
    .X(clknet_1_0__leaf_net332));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net332 (.A(clknet_0_net332),
    .X(clknet_1_1__leaf_net332));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net331 (.A(net331),
    .X(clknet_0_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net331 (.A(clknet_0_net331),
    .X(clknet_1_0__leaf_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net331 (.A(clknet_0_net331),
    .X(clknet_1_1__leaf_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net340 (.A(net340),
    .X(clknet_0_net340));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net340 (.A(clknet_0_net340),
    .X(clknet_1_0__leaf_net340));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net340 (.A(clknet_0_net340),
    .X(clknet_1_1__leaf_net340));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net801 (.A(net801),
    .X(clknet_0_net801));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net801 (.A(clknet_0_net801),
    .X(clknet_1_0__leaf_net801));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net801 (.A(clknet_0_net801),
    .X(clknet_1_1__leaf_net801));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net431 (.A(net431),
    .X(clknet_0_net431));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net431 (.A(clknet_0_net431),
    .X(clknet_1_0__leaf_net431));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net431 (.A(clknet_0_net431),
    .X(clknet_1_1__leaf_net431));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net365 (.A(net365),
    .X(clknet_0_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net365 (.A(clknet_0_net365),
    .X(clknet_1_0__leaf_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net365 (.A(clknet_0_net365),
    .X(clknet_1_1__leaf_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net460 (.A(net460),
    .X(clknet_0_net460));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net460 (.A(clknet_0_net460),
    .X(clknet_1_0__leaf_net460));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net460 (.A(clknet_0_net460),
    .X(clknet_1_1__leaf_net460));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net458 (.A(net458),
    .X(clknet_0_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net458 (.A(clknet_0_net458),
    .X(clknet_1_0__leaf_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net458 (.A(clknet_0_net458),
    .X(clknet_1_1__leaf_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net324 (.A(net324),
    .X(clknet_0_net324));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net324 (.A(clknet_0_net324),
    .X(clknet_1_0__leaf_net324));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net324 (.A(clknet_0_net324),
    .X(clknet_1_1__leaf_net324));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net328 (.A(net328),
    .X(clknet_0_net328));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net328 (.A(clknet_0_net328),
    .X(clknet_1_0__leaf_net328));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net328 (.A(clknet_0_net328),
    .X(clknet_1_1__leaf_net328));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net800 (.A(net800),
    .X(clknet_0_net800));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net800 (.A(clknet_0_net800),
    .X(clknet_1_0__leaf_net800));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net800 (.A(clknet_0_net800),
    .X(clknet_1_1__leaf_net800));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net425 (.A(net425),
    .X(clknet_0_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net425 (.A(clknet_0_net425),
    .X(clknet_1_0__leaf_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net425 (.A(clknet_0_net425),
    .X(clknet_1_1__leaf_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net439 (.A(net439),
    .X(clknet_0_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net439 (.A(clknet_0_net439),
    .X(clknet_1_0__leaf_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net439 (.A(clknet_0_net439),
    .X(clknet_1_1__leaf_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net838 (.A(net838),
    .X(clknet_0_net838));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net838 (.A(clknet_0_net838),
    .X(clknet_1_0__leaf_net838));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net838 (.A(clknet_0_net838),
    .X(clknet_1_1__leaf_net838));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net999 (.A(net999),
    .X(clknet_0_net999));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net999 (.A(clknet_0_net999),
    .X(clknet_1_0__leaf_net999));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net999 (.A(clknet_0_net999),
    .X(clknet_1_1__leaf_net999));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net493 (.A(net493),
    .X(clknet_0_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net493 (.A(clknet_0_net493),
    .X(clknet_1_0__leaf_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net493 (.A(clknet_0_net493),
    .X(clknet_1_1__leaf_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net784 (.A(net784),
    .X(clknet_0_net784));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net784 (.A(clknet_0_net784),
    .X(clknet_1_0__leaf_net784));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net784 (.A(clknet_0_net784),
    .X(clknet_1_1__leaf_net784));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net783 (.A(net783),
    .X(clknet_0_net783));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net783 (.A(clknet_0_net783),
    .X(clknet_1_0__leaf_net783));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net783 (.A(clknet_0_net783),
    .X(clknet_1_1__leaf_net783));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net396 (.A(net396),
    .X(clknet_0_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_0__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_1__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net969 (.A(net969),
    .X(clknet_0_net969));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net969 (.A(clknet_0_net969),
    .X(clknet_1_0__leaf_net969));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net969 (.A(clknet_0_net969),
    .X(clknet_1_1__leaf_net969));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net301 (.A(net301),
    .X(clknet_0_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net301 (.A(clknet_0_net301),
    .X(clknet_1_0__leaf_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net301 (.A(clknet_0_net301),
    .X(clknet_1_1__leaf_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net782 (.A(net782),
    .X(clknet_0_net782));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net782 (.A(clknet_0_net782),
    .X(clknet_1_0__leaf_net782));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net782 (.A(clknet_0_net782),
    .X(clknet_1_1__leaf_net782));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net361 (.A(net361),
    .X(clknet_0_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net361 (.A(clknet_0_net361),
    .X(clknet_1_0__leaf_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net361 (.A(clknet_0_net361),
    .X(clknet_1_1__leaf_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net976 (.A(net976),
    .X(clknet_0_net976));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net976 (.A(clknet_0_net976),
    .X(clknet_1_0__leaf_net976));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net976 (.A(clknet_0_net976),
    .X(clknet_1_1__leaf_net976));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net290 (.A(net290),
    .X(clknet_0_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net290 (.A(clknet_0_net290),
    .X(clknet_1_0__leaf_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net290 (.A(clknet_0_net290),
    .X(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net287 (.A(net287),
    .X(clknet_0_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net287 (.A(clknet_0_net287),
    .X(clknet_1_0__leaf_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net287 (.A(clknet_0_net287),
    .X(clknet_1_1__leaf_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net296 (.A(net296),
    .X(clknet_0_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net296 (.A(clknet_0_net296),
    .X(clknet_1_0__leaf_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net296 (.A(clknet_0_net296),
    .X(clknet_1_1__leaf_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net291 (.A(net291),
    .X(clknet_0_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net291 (.A(clknet_0_net291),
    .X(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net291 (.A(clknet_0_net291),
    .X(clknet_1_1__leaf_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net279 (.A(net279),
    .X(clknet_0_net279));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net279 (.A(clknet_0_net279),
    .X(clknet_1_0__leaf_net279));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net279 (.A(clknet_0_net279),
    .X(clknet_1_1__leaf_net279));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net766 (.A(net766),
    .X(clknet_0_net766));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net766 (.A(clknet_0_net766),
    .X(clknet_1_0__leaf_net766));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net766 (.A(clknet_0_net766),
    .X(clknet_1_1__leaf_net766));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net637 (.A(net637),
    .X(clknet_0_net637));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net637 (.A(clknet_0_net637),
    .X(clknet_1_0__leaf_net637));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net637 (.A(clknet_0_net637),
    .X(clknet_1_1__leaf_net637));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net990 (.A(net990),
    .X(clknet_0_net990));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net990 (.A(clknet_0_net990),
    .X(clknet_1_0__leaf_net990));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net990 (.A(clknet_0_net990),
    .X(clknet_1_1__leaf_net990));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net840 (.A(net840),
    .X(clknet_0_net840));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net840 (.A(clknet_0_net840),
    .X(clknet_1_0__leaf_net840));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net840 (.A(clknet_0_net840),
    .X(clknet_1_1__leaf_net840));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net456 (.A(net456),
    .X(clknet_0_net456));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net456 (.A(clknet_0_net456),
    .X(clknet_1_0__leaf_net456));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net456 (.A(clknet_0_net456),
    .X(clknet_1_1__leaf_net456));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net223 (.A(net223),
    .X(clknet_0_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net223 (.A(clknet_0_net223),
    .X(clknet_1_0__leaf_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net223 (.A(clknet_0_net223),
    .X(clknet_1_1__leaf_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1022 (.A(net1022),
    .X(clknet_0_net1022));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1022 (.A(clknet_0_net1022),
    .X(clknet_1_0__leaf_net1022));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1022 (.A(clknet_0_net1022),
    .X(clknet_1_1__leaf_net1022));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net325 (.A(net325),
    .X(clknet_0_net325));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net325 (.A(clknet_0_net325),
    .X(clknet_1_0__leaf_net325));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net325 (.A(clknet_0_net325),
    .X(clknet_1_1__leaf_net325));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net765 (.A(net765),
    .X(clknet_0_net765));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net765 (.A(clknet_0_net765),
    .X(clknet_1_0__leaf_net765));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net765 (.A(clknet_0_net765),
    .X(clknet_1_1__leaf_net765));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net346 (.A(net346),
    .X(clknet_0_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net346 (.A(clknet_0_net346),
    .X(clknet_1_0__leaf_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net346 (.A(clknet_0_net346),
    .X(clknet_1_1__leaf_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net996 (.A(net996),
    .X(clknet_0_net996));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net996 (.A(clknet_0_net996),
    .X(clknet_1_0__leaf_net996));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net996 (.A(clknet_0_net996),
    .X(clknet_1_1__leaf_net996));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net435 (.A(net435),
    .X(clknet_0_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net435 (.A(clknet_0_net435),
    .X(clknet_1_0__leaf_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net435 (.A(clknet_0_net435),
    .X(clknet_1_1__leaf_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net214 (.A(net214),
    .X(clknet_0_net214));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net214 (.A(clknet_0_net214),
    .X(clknet_1_0__leaf_net214));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net214 (.A(clknet_0_net214),
    .X(clknet_1_1__leaf_net214));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net202 (.A(net202),
    .X(clknet_0_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net202 (.A(clknet_0_net202),
    .X(clknet_1_0__leaf_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net202 (.A(clknet_0_net202),
    .X(clknet_1_1__leaf_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net764 (.A(net764),
    .X(clknet_0_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net764 (.A(clknet_0_net764),
    .X(clknet_1_0__leaf_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net764 (.A(clknet_0_net764),
    .X(clknet_1_1__leaf_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net232 (.A(net232),
    .X(clknet_0_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net232 (.A(clknet_0_net232),
    .X(clknet_1_0__leaf_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net232 (.A(clknet_0_net232),
    .X(clknet_1_1__leaf_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net233 (.A(net233),
    .X(clknet_0_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net233 (.A(clknet_0_net233),
    .X(clknet_1_0__leaf_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net233 (.A(clknet_0_net233),
    .X(clknet_1_1__leaf_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net745 (.A(net745),
    .X(clknet_0_net745));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net745 (.A(clknet_0_net745),
    .X(clknet_1_0__leaf_net745));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net745 (.A(clknet_0_net745),
    .X(clknet_1_1__leaf_net745));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net257 (.A(net257),
    .X(clknet_0_net257));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net257 (.A(clknet_0_net257),
    .X(clknet_1_0__leaf_net257));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net257 (.A(clknet_0_net257),
    .X(clknet_1_1__leaf_net257));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net255 (.A(net255),
    .X(clknet_0_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net255 (.A(clknet_0_net255),
    .X(clknet_1_0__leaf_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net255 (.A(net1138),
    .X(clknet_1_1__leaf_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net261 (.A(net261),
    .X(clknet_0_net261));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net261 (.A(clknet_0_net261),
    .X(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net261 (.A(clknet_0_net261),
    .X(clknet_1_1__leaf_net261));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net256 (.A(net256),
    .X(clknet_0_net256));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net256 (.A(clknet_0_net256),
    .X(clknet_1_0__leaf_net256));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net256 (.A(clknet_0_net256),
    .X(clknet_1_1__leaf_net256));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net269 (.A(net269),
    .X(clknet_0_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net269 (.A(clknet_0_net269),
    .X(clknet_1_0__leaf_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net269 (.A(clknet_0_net269),
    .X(clknet_1_1__leaf_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net744 (.A(net744),
    .X(clknet_0_net744));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net744 (.A(clknet_0_net744),
    .X(clknet_1_0__leaf_net744));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net744 (.A(clknet_0_net744),
    .X(clknet_1_1__leaf_net744));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net430 (.A(net430),
    .X(clknet_0_net430));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net430 (.A(clknet_0_net430),
    .X(clknet_1_0__leaf_net430));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net430 (.A(clknet_0_net430),
    .X(clknet_1_1__leaf_net430));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net398 (.A(net398),
    .X(clknet_0_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_0__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_1__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net400 (.A(net400),
    .X(clknet_0_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net400 (.A(clknet_0_net400),
    .X(clknet_1_0__leaf_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net400 (.A(clknet_0_net400),
    .X(clknet_1_1__leaf_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1002 (.A(net1002),
    .X(clknet_0_net1002));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1002 (.A(clknet_0_net1002),
    .X(clknet_1_0__leaf_net1002));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1002 (.A(clknet_0_net1002),
    .X(clknet_1_1__leaf_net1002));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net211 (.A(net211),
    .X(clknet_0_net211));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net211 (.A(clknet_0_net211),
    .X(clknet_1_0__leaf_net211));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net211 (.A(clknet_0_net211),
    .X(clknet_1_1__leaf_net211));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net215 (.A(net215),
    .X(clknet_0_net215));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net215 (.A(clknet_0_net215),
    .X(clknet_1_0__leaf_net215));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net215 (.A(clknet_0_net215),
    .X(clknet_1_1__leaf_net215));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net743 (.A(net743),
    .X(clknet_0_net743));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net743 (.A(clknet_0_net743),
    .X(clknet_1_0__leaf_net743));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net743 (.A(clknet_0_net743),
    .X(clknet_1_1__leaf_net743));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net503 (.A(net503),
    .X(clknet_0_net503));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net503 (.A(clknet_0_net503),
    .X(clknet_1_0__leaf_net503));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net503 (.A(clknet_0_net503),
    .X(clknet_1_1__leaf_net503));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net513 (.A(net513),
    .X(clknet_0_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net513 (.A(clknet_0_net513),
    .X(clknet_1_0__leaf_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net513 (.A(clknet_0_net513),
    .X(clknet_1_1__leaf_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net525 (.A(net525),
    .X(clknet_0_net525));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net525 (.A(clknet_0_net525),
    .X(clknet_1_0__leaf_net525));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net525 (.A(clknet_0_net525),
    .X(clknet_1_1__leaf_net525));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net519 (.A(net519),
    .X(clknet_0_net519));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net519 (.A(clknet_0_net519),
    .X(clknet_1_0__leaf_net519));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net519 (.A(clknet_0_net519),
    .X(clknet_1_1__leaf_net519));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net506 (.A(net506),
    .X(clknet_0_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net506 (.A(clknet_0_net506),
    .X(clknet_1_0__leaf_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net506 (.A(clknet_0_net506),
    .X(clknet_1_1__leaf_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net505 (.A(net505),
    .X(clknet_0_net505));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net505 (.A(clknet_0_net505),
    .X(clknet_1_0__leaf_net505));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net505 (.A(clknet_0_net505),
    .X(clknet_1_1__leaf_net505));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net504 (.A(net504),
    .X(clknet_0_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net504 (.A(clknet_0_net504),
    .X(clknet_1_0__leaf_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net504 (.A(clknet_0_net504),
    .X(clknet_1_1__leaf_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net185 (.A(net185),
    .X(clknet_0_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net185 (.A(clknet_0_net185),
    .X(clknet_1_0__leaf_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net185 (.A(clknet_0_net185),
    .X(clknet_1_1__leaf_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net193 (.A(net193),
    .X(clknet_0_net193));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net193 (.A(clknet_0_net193),
    .X(clknet_1_0__leaf_net193));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net193 (.A(clknet_0_net193),
    .X(clknet_1_1__leaf_net193));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net191 (.A(net191),
    .X(clknet_0_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net191 (.A(clknet_0_net191),
    .X(clknet_1_0__leaf_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net191 (.A(clknet_0_net191),
    .X(clknet_1_1__leaf_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net189 (.A(net189),
    .X(clknet_0_net189));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net189 (.A(clknet_0_net189),
    .X(clknet_1_0__leaf_net189));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net189 (.A(clknet_0_net189),
    .X(clknet_1_1__leaf_net189));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net197 (.A(net197),
    .X(clknet_0_net197));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net197 (.A(clknet_0_net197),
    .X(clknet_1_0__leaf_net197));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net197 (.A(clknet_0_net197),
    .X(clknet_1_1__leaf_net197));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net164 (.A(net164),
    .X(clknet_0_net164));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net164 (.A(clknet_0_net164),
    .X(clknet_1_0__leaf_net164));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net164 (.A(clknet_0_net164),
    .X(clknet_1_1__leaf_net164));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net726 (.A(net726),
    .X(clknet_0_net726));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net726 (.A(clknet_0_net726),
    .X(clknet_1_0__leaf_net726));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net726 (.A(clknet_0_net726),
    .X(clknet_1_1__leaf_net726));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net725 (.A(net725),
    .X(clknet_0_net725));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net725 (.A(clknet_0_net725),
    .X(clknet_1_0__leaf_net725));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net725 (.A(clknet_0_net725),
    .X(clknet_1_1__leaf_net725));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net112 (.A(net112),
    .X(clknet_0_net112));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net112 (.A(clknet_0_net112),
    .X(clknet_1_0__leaf_net112));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net112 (.A(clknet_0_net112),
    .X(clknet_1_1__leaf_net112));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net102 (.A(net102),
    .X(clknet_0_net102));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net102 (.A(clknet_0_net102),
    .X(clknet_1_0__leaf_net102));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net102 (.A(clknet_0_net102),
    .X(clknet_1_1__leaf_net102));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net987 (.A(net987),
    .X(clknet_0_net987));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net987 (.A(clknet_0_net987),
    .X(clknet_1_0__leaf_net987));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net987 (.A(clknet_0_net987),
    .X(clknet_1_1__leaf_net987));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net117 (.A(net117),
    .X(clknet_0_net117));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net117 (.A(clknet_0_net117),
    .X(clknet_1_0__leaf_net117));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net117 (.A(clknet_0_net117),
    .X(clknet_1_1__leaf_net117));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net113 (.A(net113),
    .X(clknet_0_net113));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net113 (.A(clknet_0_net113),
    .X(clknet_1_0__leaf_net113));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net113 (.A(clknet_0_net113),
    .X(clknet_1_1__leaf_net113));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net100 (.A(net100),
    .X(clknet_0_net100));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net100 (.A(clknet_0_net100),
    .X(clknet_1_0__leaf_net100));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net100 (.A(clknet_0_net100),
    .X(clknet_1_1__leaf_net100));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net104 (.A(net104),
    .X(clknet_0_net104));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net104 (.A(clknet_0_net104),
    .X(clknet_1_0__leaf_net104));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net104 (.A(clknet_0_net104),
    .X(clknet_1_1__leaf_net104));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net206 (.A(net206),
    .X(clknet_0_net206));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net206 (.A(clknet_0_net206),
    .X(clknet_1_0__leaf_net206));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net206 (.A(clknet_0_net206),
    .X(clknet_1_1__leaf_net206));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net103 (.A(net103),
    .X(clknet_0_net103));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net103 (.A(clknet_0_net103),
    .X(clknet_1_0__leaf_net103));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net103 (.A(clknet_0_net103),
    .X(clknet_1_1__leaf_net103));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net724 (.A(net724),
    .X(clknet_0_net724));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net724 (.A(clknet_0_net724),
    .X(clknet_1_0__leaf_net724));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net724 (.A(clknet_0_net724),
    .X(clknet_1_1__leaf_net724));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net705 (.A(net705),
    .X(clknet_0_net705));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net705 (.A(clknet_0_net705),
    .X(clknet_1_0__leaf_net705));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net705 (.A(clknet_0_net705),
    .X(clknet_1_1__leaf_net705));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net181 (.A(net181),
    .X(clknet_0_net181));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net181 (.A(clknet_0_net181),
    .X(clknet_1_0__leaf_net181));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net181 (.A(clknet_0_net181),
    .X(clknet_1_1__leaf_net181));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net404 (.A(net404),
    .X(clknet_0_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net404 (.A(clknet_0_net404),
    .X(clknet_1_0__leaf_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net404 (.A(clknet_0_net404),
    .X(clknet_1_1__leaf_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net183 (.A(net183),
    .X(clknet_0_net183));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net183 (.A(clknet_0_net183),
    .X(clknet_1_0__leaf_net183));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net183 (.A(clknet_0_net183),
    .X(clknet_1_1__leaf_net183));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net88 (.A(net88),
    .X(clknet_0_net88));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net88 (.A(clknet_0_net88),
    .X(clknet_1_0__leaf_net88));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net88 (.A(clknet_0_net88),
    .X(clknet_1_1__leaf_net88));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net635 (.A(net635),
    .X(clknet_0_net635));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net635 (.A(clknet_0_net635),
    .X(clknet_1_0__leaf_net635));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net635 (.A(clknet_0_net635),
    .X(clknet_1_1__leaf_net635));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1003 (.A(net1003),
    .X(clknet_0_net1003));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1003 (.A(clknet_0_net1003),
    .X(clknet_1_0__leaf_net1003));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1003 (.A(clknet_0_net1003),
    .X(clknet_1_1__leaf_net1003));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net82 (.A(net82),
    .X(clknet_0_net82));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net82 (.A(clknet_0_net82),
    .X(clknet_1_0__leaf_net82));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net82 (.A(clknet_0_net82),
    .X(clknet_1_1__leaf_net82));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net83 (.A(net83),
    .X(clknet_0_net83));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net83 (.A(clknet_0_net83),
    .X(clknet_1_0__leaf_net83));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net83 (.A(clknet_0_net83),
    .X(clknet_1_1__leaf_net83));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net979 (.A(net979),
    .X(clknet_0_net979));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net979 (.A(clknet_0_net979),
    .X(clknet_1_0__leaf_net979));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net979 (.A(clknet_0_net979),
    .X(clknet_1_1__leaf_net979));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net704 (.A(net704),
    .X(clknet_0_net704));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net704 (.A(clknet_0_net704),
    .X(clknet_1_0__leaf_net704));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net704 (.A(clknet_0_net704),
    .X(clknet_1_1__leaf_net704));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net217 (.A(net217),
    .X(clknet_0_net217));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net217 (.A(clknet_0_net217),
    .X(clknet_1_0__leaf_net217));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net217 (.A(clknet_0_net217),
    .X(clknet_1_1__leaf_net217));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net241 (.A(net241),
    .X(clknet_0_net241));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net241 (.A(clknet_0_net241),
    .X(clknet_1_0__leaf_net241));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net241 (.A(clknet_0_net241),
    .X(clknet_1_1__leaf_net241));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net225 (.A(net225),
    .X(clknet_0_net225));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net225 (.A(clknet_0_net225),
    .X(clknet_1_0__leaf_net225));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net225 (.A(clknet_0_net225),
    .X(clknet_1_1__leaf_net225));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net703 (.A(net703),
    .X(clknet_0_net703));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net703 (.A(clknet_0_net703),
    .X(clknet_1_0__leaf_net703));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net703 (.A(clknet_0_net703),
    .X(clknet_1_1__leaf_net703));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net277 (.A(net277),
    .X(clknet_0_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net277 (.A(clknet_0_net277),
    .X(clknet_1_0__leaf_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net277 (.A(clknet_0_net277),
    .X(clknet_1_1__leaf_net277));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net627),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net1128),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net1128),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net627),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net1131),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net627),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net1174),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net1134),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net1134),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net746),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(clknet_0_net255),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net855),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net755),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net761),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net708),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net781),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net700),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net756),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net600),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net610),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net697),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net1036),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net848),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net1046),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net20),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net842),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net847),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net259),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net495),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net147),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net148),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net830),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net371),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net683),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net1083),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net780),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net152),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net28),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net988),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net699),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net266),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net1047),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net849),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net751),
    .X(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in62));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in63));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in64));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(in65));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(in66));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(in67));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(in68));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(in69));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(in70));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(in71));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(in72));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(in73));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(in74));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(in75));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(in76));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(in77));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(in78));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(in79));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(in80));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(in81));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(in82));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(in83));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(in84));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(in85));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(in86));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(in87));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(in88));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(in89));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(in90));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(in91));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(in92));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(in93));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(in94));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(in95));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(in96));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(in97));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(in98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(in99));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net100_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_X (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_D (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_SCD (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_RESET_B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_SCE (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_X (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A3 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_SCE (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_SCD (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_Q_N (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A0 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_Q (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A3 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_Q_N (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_D (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_Q (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_S0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_Q (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_S1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_Q_N (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A0 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_Q (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S0 (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S0 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A0 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_X (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold30_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A3 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A3 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_Q_N (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold31_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_Q (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A0 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A0 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A0 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_X (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold37_A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_Q (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_D (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_SCD (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_X (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A3 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_SCD (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_Q_N (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A0 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A0 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A0 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_Q (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A0 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A3 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A3 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A3 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_X (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A0 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_S0 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_X (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A3 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A3 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_Q_N (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A0 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A0 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_Q (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A0 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A0 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A0 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_X (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A3 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A3 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A3 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_Q_N (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A0 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A0 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_Q (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_X (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A0 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A4 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_RESET_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A0 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_X (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A0 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A3 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_D (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A0 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A3 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A4 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_X (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_X (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A0 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_Q (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A3 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_D (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_D (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_SET_B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_X (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A3 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A3 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_Q_N (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A0 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A0 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_D (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_Q (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A3 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_X (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_SCE (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A0 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_D (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A3 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_RESET_B (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_D (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_X (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net261_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_X (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A3 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_SCD (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A3 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_SCD (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_Q_N (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A0 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_S0 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_Q (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A3 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A3 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_Q_N (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A0 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A0 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_Q (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A0 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A3 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A0 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_Q (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A0 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_D (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A0 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_RESET_B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A0 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_X (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_X (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A0 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A3 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_RESET_B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A3 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S0 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_Q_N (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A0 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A0 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A0 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_Q (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold38_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_SCD (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_S0 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_Q_N (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A0 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A0 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A0 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_Q (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A3 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S0 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A2 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A2 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_Q (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A0 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A0 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_Q (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A0 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_Q (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net291_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_X (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A3 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_X (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A0 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A0 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A3 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A3 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_X (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A0 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A3 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A3 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_X (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_X (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A3 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_S0 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S0 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_Q_N (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_Q (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S0 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A3 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_RESET_B (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A3 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_Q_N (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A0 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A2 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_D (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A0 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_Q (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_X (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A0 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A0 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_Q_N (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_RESET_B (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_S0 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A2 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_Q_N (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A0 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A0 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_Q (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A0 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A3 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A0 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A0 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_D (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_X (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_S0 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_SCD (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A4 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A3 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A3 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A3 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_SCE (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_S0 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_Q_N (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A3 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_SCD (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_SCD (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A3 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_SCD (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_Q_N (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net390_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_X (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A2 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A1 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A1 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A2 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_X (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A3 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A3 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_Q (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A1 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_X (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap221_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A4 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_S0 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_Q_N (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_Q (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_B (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_X (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A3 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A0 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_SCD (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_X (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A0 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A3 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_S0 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_S1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A4 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_SET_B (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_Q_N (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A2 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_X (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_S0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_Q (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A0 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_S0 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A3 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_D (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_S0 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_SCE (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_SCD (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_X (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A2 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A0 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A2 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_Q_N (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net505_A (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_X (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A2 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A2 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_X (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_S0 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A3 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_Q_N (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge885_D (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_X (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_X (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_X (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_B (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_X (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_S0 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A3 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_S0 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A3 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A4 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A3 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_Q_N (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_Q (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap218_A (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_Q (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_S1 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A3 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S0 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B1 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold19_A (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_Q (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_SCE (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A2 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_S0 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A4 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_S0 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_SCE (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_B (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_Y (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_Q (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A4 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_S1 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S0 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A3 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A3 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_Q (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_S0 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_S0 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold20_A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_Q_N (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_S0 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A3 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_S0 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A4 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_S1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_S0 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_Q (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A4 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_SCE (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_SCD (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_S1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A2 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A2 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_S0 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_S1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_S0 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_S0 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_Q (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A2 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A3 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_SCE (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_S0 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_SCE (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_Q (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_S1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A3 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_S0 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S0 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_S1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A3 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A4 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_Q (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A3 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A1 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A1 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S0 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A2 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A2 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S0 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_S0 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A3 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_S1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_SCE (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_S0 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_S0 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A3 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_Q (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A3 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A3 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A3 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A3 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net635_A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_GCLK (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A0 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_X (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A3 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A3 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A2 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S0 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A2 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_Q (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A3 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A3 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_Q_N (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A2 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge864_Q (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A2 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_S1 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A3 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_Q (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A3 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S1 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A3 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A2 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_Q (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A3 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S1 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_S1 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A2 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S0 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_S0 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_D (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_X (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_Q (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A3 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge885_Q (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A3 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A3 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A3 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge886_Q (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_S0 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_S0 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_S0 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S0 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S0 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_SCE (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge888_Q_N (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S0 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_Q_N (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A2 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B1 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A3 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_S1 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_S1 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_SET_B (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold21_A (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_Q (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A3 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_S0 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_SCE (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_S1 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold40_A (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_Q (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_S0 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A4 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S0 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_S1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold17_A (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_Q (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_S0 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A2 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_S0 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A4 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A4 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_SET_B (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_SET_B (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_Q (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_Q (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net703_A (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_GCLK (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net704_A (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_GCLK (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_Q_N (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A3 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A3 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_B1 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S1 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_Q (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A2 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A2 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_S1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_Q_N (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S0 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_S0 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_S0 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_S1 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_Q (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S0 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_S0 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S1 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_S0 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_Q (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A3 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S0 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A3 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A2 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_S0 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_S1 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A2 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A4 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_B1 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_Q (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_S0 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A2 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A3 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S0 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_S1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_S1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_S1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_Q (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A3 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S0 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S0 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_S1 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A3 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_S1 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S1 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S1 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B1 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap212_A (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_Q (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A3 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A3 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S0 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_S1 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_S1 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap211_A (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_s905_Q (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_S0 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S1 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_Q_N (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S0 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_Q (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S0 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A3 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A2 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_Q_N (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S0 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_S0 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_S0 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A3 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_Q (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A2 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A3 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_S1 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_s908_Q (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S0 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A3 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S0 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S0 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_S1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_Q (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A3 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S0 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A3 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_S0 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_S0 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_Q (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S0 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_X (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_Q (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_Q (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_S0 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A2 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_S0 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_S1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_S1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_Q (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A2 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S0 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S1 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_S1 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_S1 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_S1 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_S1 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_s921_Q (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A1 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S0 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A3 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S0 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_S0 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_Q_N (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A2 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_S0 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A3 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_X (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_s924_Q (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A3 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_S1 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_S1 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_S1 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_Q (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S1 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S1 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S0 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A3 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S1 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net745_A (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_s929_GCLK (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_Q (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_SET_B (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S0 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A3 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_Q_N (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S0 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A3 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_S0 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_Q (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S0 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_s933_Q (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_S1 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S0 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A3 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_S0 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_S0 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_S1 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_B1 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_S1 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_S0 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_S1 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_Q (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S0 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_S0 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_S0 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_S1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_s935_Q (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A1 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_S1 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S0 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A3 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S0 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold18_A (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_Q (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_S0 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_S1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S0 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_S1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_S1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_s939_Q_N (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A3 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A3 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_S1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_S1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_S1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A3 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_X (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_s939_Q (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_S0 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S0 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A3 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_S0 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_S1 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold14_A (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_s940_Q (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S0 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S0 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_S1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_S1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_s941_Q (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A2 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S0 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A3 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S0 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_S0 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S0 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_s942_Q (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S0 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S0 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_S0 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_s946_Q_N (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S0 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A3 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_s950_Q (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A3 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S0 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S0 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_S0 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_s951_Q (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S0 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S0 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A3 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S0 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_S1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_SCE (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_X (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold36_A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_s957_Q (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A3 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A2 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_S1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A4 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_S1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_S1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net783_A (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_s960_GCLK (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_s962_Q (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_S0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A3 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_S1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_s963_Q_N (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_S1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_s964_Q (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_S0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_S1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_S0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A3 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_s967_Q (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A3 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_S1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_S1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_s968_Q (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_SET_B (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A3 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_s971_Q_N (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A3 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_S1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A3 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_s971_Q (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S0 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S0 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_s974_Q (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S0 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_s982_Q (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_B1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_s988_Q (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A3 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S0 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_S1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_s989_Q (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A3 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A3 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_S0 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A4 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_B1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_s990_Q (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A3 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A3 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_S0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A4 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_s996_Q (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_S1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_s997_Q (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_S1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_s999_Q (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_S1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_s1003_Q (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A3 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold23_A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_s1015_Q (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A3 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_S0 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_SET_B (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_s1018_Q_N (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_S1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_s1018_Q (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_S0 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_s1019_Q (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S1 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_S0 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_s1021_Q (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S0 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_S1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_S1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_S1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_S1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_S1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_s1022_Q (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_S0 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_S1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S0 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_A (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A3 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A2 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A0 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A3 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A3 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A0 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A2 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_RESET_B (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_D (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A2 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A2 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A2 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A3 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S0 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_A (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_A (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A0 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A2 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A2 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A0 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_SCD (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A3 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A0 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A3 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A3 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_S0 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A3 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A0 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A2 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A3 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A2 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_A (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_A (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A0 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A0 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_S1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A2 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A2 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A3 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A3 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A2 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_S1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A2 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_D (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_S0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_B1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A0 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A2 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A0 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A3 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A3 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A3 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A2 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A0 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A2 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A2 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A0 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A2 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A0 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_D (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A0 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A4 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_S1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_S1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A3 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A0 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A2 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A0 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A0 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A0 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A0 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A3 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A0 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A0 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A3 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A4 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A2 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A3 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A0 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A3 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A3 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_S1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_S0 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A0 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_SCD (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_A3 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A0 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A2 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A2 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_RESET_B (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_X (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A0 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A2 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A2 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_S0 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_S0 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_D (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_S0 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A0 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A0 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A2 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_S0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A1 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A0 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A0 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A2 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A2 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A1 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A1 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A0 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A0 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A4 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A0 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A3 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A3 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_S0 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_A (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A2 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_D (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A1 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A1 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A3 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A2 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A2 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A2 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A0 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A2 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A1 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A3 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A0 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_S0 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A0 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S0 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A2 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A3 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A1 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A2 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A3 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A2 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A1 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_S1 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A0 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A3 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_S0 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_S1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_X (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_S0 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A3 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A4 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_SET_B (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_S1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A2 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S0 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A0 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A3 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A2 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_S0 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_B1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_B1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A3 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_A (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A2 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A1 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A0 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A3 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A2 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A3 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_X (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A0 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A0 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A4 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_S0 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S0 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A3 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A2 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A2 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A0 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A0 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A0 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A2 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A2 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A2 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_X (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A0 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S0 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A3 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_X (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A0 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A3 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A3 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_X (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_S1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_SCD (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A3 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_X (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_X (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_B1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_A0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_S1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_S1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_X (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A0 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A2 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_X (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A0 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A0 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A0 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S0 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_X (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A0 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A0 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A3 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_X (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A2 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_X (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A0 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S0 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A0 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A0 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_X (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A2 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A0 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A0 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A2 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A3 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_X (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_X (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A0 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A0 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_X (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A0 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A3 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A3 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A3 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_X (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A2 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_X (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A0 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A0 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_SCD (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A2 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_X (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A2 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A0 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A0 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A3 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A2 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_S0 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_X (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_X (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A3 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A3 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A3 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_S0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_S0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_X (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_S0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_X (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A0 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_X (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net969_A (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_X (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_Q (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_Q (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_S0 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S0 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_RESET_B (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A3 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A3 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_S0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_SCD (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_Q (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_s979_Q (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_S1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A4 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_s963_Q (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A3 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A3 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A2 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_S1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_B1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net979_A (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_X (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_Q (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge889_Q_N (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A2 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap222_A (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A0 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_Q (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A2 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S0 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A3 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A0 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_X (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_s1006_Q (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A3 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net990_A (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_X (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_Q (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net992_A (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_X (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_s1011_Q (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_S1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net996_A (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_X (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_output130_A (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_Q (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A3 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_S1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net999_A (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_GCLK (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_output134_A (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_Q (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A3 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net1002_A (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_X (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net1003_A (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_X (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_output137_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_Q (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A3 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A3 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_S0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_output139_A (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_Q (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_output140_A (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_s949_Q (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_S0 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_output141_A (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A3 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_X (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_A (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A2 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_Q (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_output144_A (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_s969_Q (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S0 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_output145_A (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_Q (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_SCE (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_output147_A (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge847_Q (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A3 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A3 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A3 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_output148_A (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_s973_Q (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_S0 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_output149_A (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A3 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A3 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_Q (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_output154_A (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A2 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_X (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_output156_A (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_Q (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A3 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_S0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_S0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_S0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_S1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_output161_A (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_S0 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_Q (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_output168_A (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A0 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_X (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold22_A (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_output169_A (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_Q (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A3 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A3 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_S0 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_output172_A (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A1 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_output173_A (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_Q (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_S0 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S0 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_output175_A (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_S0 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A3 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S0 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A3 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_X (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_X (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A0 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_RESET_B (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A2 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_SCE (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_SET_B (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_D (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_X (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S0 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_SCD (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_SCE (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_RESET_B (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A3 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A2 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A3 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A1 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A1 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A3 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_X (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A3 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_SCE (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_S0 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A0 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_SCD (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_SCE (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A1 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_SET_B (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_SCE (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_RESET_B (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_X (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A1 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A1 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_RESET_B (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A0 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A2 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_X (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A1 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_SCD (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A1 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A3 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A3 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A2 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A1 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S0 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A3 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A4 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_X (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S0 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A2 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S0 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_S1 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A2 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A2 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A3 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A2 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A2 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A0 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_X (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A3 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A1 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_SCE (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A0 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A2 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A1 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_SCD (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_SCD (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A0 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_X (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A2 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A2 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A3 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_D (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_SET_B (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A1 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_SCE (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_SET_B (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_X (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A0 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A1 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A0 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A2 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_D (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A2 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_RESET_B (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_D (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A3 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_X (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A2 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_SCD (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_SCE (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A4 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_RESET_B (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_D (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A2 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A0 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A3 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_SCD (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_X (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_S1 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A0 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_X (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A1 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A0 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_RESET_B (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A3 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A0 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A1 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A3 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A2 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_SCE (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_X (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A2 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A1 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A3 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A2 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A1 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_X (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A2 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A2 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A2 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A1 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A2 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A1 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A2 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_S1 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A2 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A0 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_X (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A2 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A3 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A3 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A3 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_X (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A0 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S0 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A3 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_S1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A0 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_X (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S0 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A1 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A0 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A2 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A3 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A3 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_X (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A1 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A1 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A1 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A2 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_X (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A0 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A0 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A3 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_RESET_B (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_RESET_B (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A2 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A3 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B1 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_X (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A2 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A3 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A3 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A2 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A2 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A2 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A3 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_S1 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A1 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A3 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_X (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A2 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A3 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A1 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A2 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A0 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A4 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_S0 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A3 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_SCE (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A3 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_X (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A0 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A2 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A2 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A3 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S0 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A3 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_X (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A0 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A1 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_SCD (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A3 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A1 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A1 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A2 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_SET_B (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A1 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B1 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_X (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A2 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_D (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_RESET_B (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A2 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A4 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B1 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A0 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A3 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S0 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A2 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_X (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S0 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S0 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S0 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A3 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_S0 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S0 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_S0 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire209_X (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S1 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S0 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_S0 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A3 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S1 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S0 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_X (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_S0 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S0 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A3 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_S1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S0 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_S0 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_S1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_S1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap211_X (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A3 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A3 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap212_X (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S0 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_S1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_X (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A3 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A3 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_B1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S0 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_S1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_S1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_S1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_SET_B (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A3 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_X (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S0 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A3 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_S0 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_S0 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_X (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_S1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A3 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_SET_B (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_SCE (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A3 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_B1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_S0 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S0 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold35_A (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_X (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_S1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_S1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_S1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap217_X (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_S0 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S0 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S1 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S1 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S1 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S0 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S0 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap218_X (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_S0 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A3 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_S1 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A3 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_S0 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A3 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_X (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_S0 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_SCD (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A2 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A2 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A3 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A2 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_S0 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_S0 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A4 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_X (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A1 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A0 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A2 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_SET_B (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A2 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A2 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_RESET_B (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A2 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A2 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap221_X (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A2 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A2 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A3 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap222_X (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A3 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A1 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A0 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_X (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A3 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_S0 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A4 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_RESET_B (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_S0 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_SCD (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A3 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B1 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_SCE (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_S0 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_X (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_RESET_B (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A3 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A0 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A2 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A3 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A4 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_RESET_B (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_X (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A2 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_S0 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A2 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A0 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A3 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_SCD (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A3 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_X (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_SCE (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A1 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A3 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A2 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_S0 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_S1 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_SCD (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A1 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A3 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A2 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_X (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_B1 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_SCD (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_RESET_B (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B1 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A4 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_D (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_RESET_B (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A1 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A1 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A4 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_X (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B1 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_SCD (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A1 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_RESET_B (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A4 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_RESET_B (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A0 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A2 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A2 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A4 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_X (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A0 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A3 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_S1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_A4 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_X (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A2 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A3 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_S0 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A1 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A2 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A1 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_RESET_B (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A2 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_X (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A2 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A2 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A4 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B1 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A3 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_X (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S0 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A1 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A2 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A2 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A3 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_B1 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_S0 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_S0 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_D (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A1 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_X (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A2 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A1 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A2 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_SCD (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A1 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_SCE (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S0 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A0 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_SCD (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A1 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_X (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A1 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A1 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_X (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A1 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A0 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_SCD (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A1 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A3 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_S0 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A1 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_D (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A3 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_X (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A1 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A0 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_SET_B (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A2 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S1 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_X (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A2 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_RESET_B (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A3 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A3 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A1 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A0 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S1 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A2 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A3 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_S1 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_X (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S0 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S0 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A2 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_X (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A0 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A3 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A3 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A0 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A4 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A2 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_D (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A3 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_X (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A3 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_S1 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A0 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_SCE (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A1 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A1 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A2 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A0 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A1 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A3 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_X (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A3 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A3 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A0 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A1 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_SCE (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A0 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_SCD (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A1 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_D (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A3 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_X (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A0 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A1 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A3 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S0 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A1 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A0 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A3 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A2 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A2 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_X (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S0 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S0 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A1 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A0 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A2 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A2 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A1 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A1 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A1 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_X (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A4 (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S0 (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_SCE (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A3 (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A2 (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A4 (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_RESET_B (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B1 (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A4 (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B1 (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_X (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A2 (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S0 (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A2 (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A2 (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B1 (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B1 (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_X (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A0 (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_S1 (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_B1 (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_D (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_A3 (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_S0 (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_B1 (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_S1 (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A3 (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A3 (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_X (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_A (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A2 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A3 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A0 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_X (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A2 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A2 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A3 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A2 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A3 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_S0 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A3 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_S0 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_SCE (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_SET_B (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_X (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A3 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A2 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S0 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_S0 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A3 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_X (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A1 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A0 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_SCD (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A1 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_S1 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A3 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A1 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A1 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A2 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B1 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_X (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A2 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A3 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_SET_B (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A1 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A4 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A1 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A3 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_S1 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_S0 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A3 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_X (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A1 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A1 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S0 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A0 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_X (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A1 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A2 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A1 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_S0 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A3 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A1 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A2 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A2 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A3 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A3 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_X (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A1 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A2 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A3 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A1 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_S0 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A2 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A1 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A1 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A3 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A3 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_X (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A1 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_S0 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A0 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A1 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A0 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_SCD (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A0 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_S1 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_S0 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B1 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_X (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A0 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A1 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_D (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A1 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_S0 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A1 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A2 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A2 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A1 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_SCD (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_X (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A4 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A1 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A3 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A1 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A0 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A1 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_S0 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A2 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A1 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A3 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_X (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A0 (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A3 (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A3 (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_S1 (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A3 (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A0 (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A1 (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_D (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A4 (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A2 (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_X (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A1 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A2 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S0 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A3 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A2 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S0 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A0 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_S0 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A3 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A3 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_X (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A3 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A2 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A2 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_D (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A1 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A0 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A3 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_B1 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A3 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_X (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s1000_GATE (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_X (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_X (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_X (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net818_A (.DIODE(clknet_0_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net818_A (.DIODE(clknet_0_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net818_X (.DIODE(clknet_0_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_B1 (.DIODE(clknet_1_0__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_S1 (.DIODE(clknet_1_0__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_B1 (.DIODE(clknet_1_0__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_B1 (.DIODE(clknet_1_0__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_S0 (.DIODE(clknet_1_0__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_S1 (.DIODE(clknet_1_0__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_S1 (.DIODE(clknet_1_0__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_B1 (.DIODE(clknet_1_0__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_S0 (.DIODE(clknet_1_0__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net818_X (.DIODE(clknet_1_0__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S1 (.DIODE(clknet_1_1__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S0 (.DIODE(clknet_1_1__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S0 (.DIODE(clknet_1_1__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S0 (.DIODE(clknet_1_1__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(clknet_1_1__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S0 (.DIODE(clknet_1_1__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(clknet_1_1__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net818_X (.DIODE(clknet_1_1__leaf_net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A3 (.DIODE(clknet_1_0__leaf_net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A0 (.DIODE(clknet_1_0__leaf_net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net393_X (.DIODE(clknet_1_0__leaf_net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S1 (.DIODE(clknet_1_0__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_SET_B (.DIODE(clknet_1_0__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(clknet_1_0__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S0 (.DIODE(clknet_1_0__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net801_X (.DIODE(clknet_1_0__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(clknet_1_1__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S1 (.DIODE(clknet_1_1__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A3 (.DIODE(clknet_1_1__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net801_X (.DIODE(clknet_1_1__leaf_net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A1 (.DIODE(clknet_1_0__leaf_net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(clknet_1_0__leaf_net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net324_X (.DIODE(clknet_1_0__leaf_net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(clknet_1_0__leaf_net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(clknet_1_0__leaf_net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A3 (.DIODE(clknet_1_0__leaf_net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net999_X (.DIODE(clknet_1_0__leaf_net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_SET_B (.DIODE(clknet_1_1__leaf_net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_SET_B (.DIODE(clknet_1_1__leaf_net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_S1 (.DIODE(clknet_1_1__leaf_net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(clknet_1_1__leaf_net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net999_X (.DIODE(clknet_1_1__leaf_net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S0 (.DIODE(clknet_1_1__leaf_net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(clknet_1_1__leaf_net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_S0 (.DIODE(clknet_1_1__leaf_net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net783_X (.DIODE(clknet_1_1__leaf_net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_S1 (.DIODE(clknet_1_1__leaf_net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_S1 (.DIODE(clknet_1_1__leaf_net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S0 (.DIODE(clknet_1_1__leaf_net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net782_X (.DIODE(clknet_1_1__leaf_net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(clknet_1_1__leaf_net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A3 (.DIODE(clknet_1_1__leaf_net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A0 (.DIODE(clknet_1_1__leaf_net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net291_X (.DIODE(clknet_1_1__leaf_net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A1 (.DIODE(clknet_1_0__leaf_net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A1 (.DIODE(clknet_1_0__leaf_net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A3 (.DIODE(clknet_1_0__leaf_net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(clknet_1_0__leaf_net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(clknet_1_0__leaf_net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(clknet_1_0__leaf_net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net990_X (.DIODE(clknet_1_0__leaf_net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A3 (.DIODE(clknet_1_1__leaf_net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(clknet_1_1__leaf_net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S0 (.DIODE(clknet_1_1__leaf_net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(clknet_1_1__leaf_net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net990_X (.DIODE(clknet_1_1__leaf_net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A2 (.DIODE(clknet_1_0__leaf_net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S0 (.DIODE(clknet_1_0__leaf_net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A3 (.DIODE(clknet_1_0__leaf_net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A2 (.DIODE(clknet_1_0__leaf_net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A3 (.DIODE(clknet_1_0__leaf_net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net1022_X (.DIODE(clknet_1_0__leaf_net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(clknet_1_1__leaf_net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_output155_A (.DIODE(clknet_1_1__leaf_net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net1022_X (.DIODE(clknet_1_1__leaf_net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A0 (.DIODE(clknet_1_0__leaf_net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A2 (.DIODE(clknet_1_0__leaf_net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_S0 (.DIODE(clknet_1_0__leaf_net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A1 (.DIODE(clknet_1_0__leaf_net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net996_X (.DIODE(clknet_1_0__leaf_net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S0 (.DIODE(clknet_1_1__leaf_net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A1 (.DIODE(clknet_1_1__leaf_net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_output129_A (.DIODE(clknet_1_1__leaf_net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net996_X (.DIODE(clknet_1_1__leaf_net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A1 (.DIODE(clknet_1_1__leaf_net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A1 (.DIODE(clknet_1_1__leaf_net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_D (.DIODE(clknet_1_1__leaf_net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A1 (.DIODE(clknet_1_1__leaf_net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net202_X (.DIODE(clknet_1_1__leaf_net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_S1 (.DIODE(clknet_1_1__leaf_net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_S1 (.DIODE(clknet_1_1__leaf_net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S1 (.DIODE(clknet_1_1__leaf_net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net764_X (.DIODE(clknet_1_1__leaf_net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(clknet_1_1__leaf_net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A3 (.DIODE(clknet_1_1__leaf_net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_S0 (.DIODE(clknet_1_1__leaf_net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S1 (.DIODE(clknet_1_1__leaf_net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net745_X (.DIODE(clknet_1_1__leaf_net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A1 (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A1 (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A1 (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A1 (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A1 (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net255_X (.DIODE(clknet_1_0__leaf_net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net261_A (.DIODE(clknet_0_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net261_A (.DIODE(clknet_0_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net261_X (.DIODE(clknet_0_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_SET_B (.DIODE(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A1 (.DIODE(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_D (.DIODE(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A3 (.DIODE(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_SCD (.DIODE(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_D (.DIODE(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A1 (.DIODE(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A2 (.DIODE(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net261_X (.DIODE(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A2 (.DIODE(clknet_1_1__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(clknet_1_1__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S0 (.DIODE(clknet_1_1__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(clknet_1_1__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(clknet_1_1__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net261_X (.DIODE(clknet_1_1__leaf_net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S0 (.DIODE(clknet_1_0__leaf_net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A3 (.DIODE(clknet_1_0__leaf_net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net744_X (.DIODE(clknet_1_0__leaf_net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_RESET_B (.DIODE(clknet_1_0__leaf_net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(clknet_1_0__leaf_net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(clknet_1_0__leaf_net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net1002_X (.DIODE(clknet_1_0__leaf_net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net743_A (.DIODE(clknet_0_net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net743_A (.DIODE(clknet_0_net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net743_X (.DIODE(clknet_0_net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_S1 (.DIODE(clknet_1_0__leaf_net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S1 (.DIODE(clknet_1_0__leaf_net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S1 (.DIODE(clknet_1_0__leaf_net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B1 (.DIODE(clknet_1_0__leaf_net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_S1 (.DIODE(clknet_1_0__leaf_net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_S0 (.DIODE(clknet_1_0__leaf_net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_S1 (.DIODE(clknet_1_0__leaf_net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net743_X (.DIODE(clknet_1_0__leaf_net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A3 (.DIODE(clknet_1_1__leaf_net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A3 (.DIODE(clknet_1_1__leaf_net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_S1 (.DIODE(clknet_1_1__leaf_net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_S1 (.DIODE(clknet_1_1__leaf_net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S0 (.DIODE(clknet_1_1__leaf_net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S0 (.DIODE(clknet_1_1__leaf_net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_S0 (.DIODE(clknet_1_1__leaf_net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net743_X (.DIODE(clknet_1_1__leaf_net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A1 (.DIODE(clknet_1_1__leaf_net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A0 (.DIODE(clknet_1_1__leaf_net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A2 (.DIODE(clknet_1_1__leaf_net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A2 (.DIODE(clknet_1_1__leaf_net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net197_X (.DIODE(clknet_1_1__leaf_net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A3 (.DIODE(clknet_1_1__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A0 (.DIODE(clknet_1_1__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A1 (.DIODE(clknet_1_1__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A0 (.DIODE(clknet_1_1__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net100_X (.DIODE(clknet_1_1__leaf_net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S1 (.DIODE(clknet_1_0__leaf_net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S0 (.DIODE(clknet_1_0__leaf_net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_S0 (.DIODE(clknet_1_0__leaf_net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_S1 (.DIODE(clknet_1_0__leaf_net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S0 (.DIODE(clknet_1_0__leaf_net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net705_X (.DIODE(clknet_1_0__leaf_net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A0 (.DIODE(clknet_1_0__leaf_net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A0 (.DIODE(clknet_1_0__leaf_net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net181_X (.DIODE(clknet_1_0__leaf_net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A2 (.DIODE(clknet_1_0__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A2 (.DIODE(clknet_1_0__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_S0 (.DIODE(clknet_1_0__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A0 (.DIODE(clknet_1_0__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A3 (.DIODE(clknet_1_0__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A1 (.DIODE(clknet_1_0__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A1 (.DIODE(clknet_1_0__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A1 (.DIODE(clknet_1_0__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(clknet_1_0__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A2 (.DIODE(clknet_1_0__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A3 (.DIODE(clknet_1_0__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_S0 (.DIODE(clknet_1_0__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A3 (.DIODE(clknet_1_0__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A1 (.DIODE(clknet_1_0__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net88_X (.DIODE(clknet_1_0__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A3 (.DIODE(clknet_1_1__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A2 (.DIODE(clknet_1_1__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A3 (.DIODE(clknet_1_1__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A0 (.DIODE(clknet_1_1__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A2 (.DIODE(clknet_1_1__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A2 (.DIODE(clknet_1_1__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A0 (.DIODE(clknet_1_1__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A2 (.DIODE(clknet_1_1__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A1 (.DIODE(clknet_1_1__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net88_X (.DIODE(clknet_1_1__leaf_net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net635_A (.DIODE(clknet_0_net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net635_A (.DIODE(clknet_0_net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net635_X (.DIODE(clknet_0_net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_S1 (.DIODE(clknet_1_0__leaf_net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_S0 (.DIODE(clknet_1_0__leaf_net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A1 (.DIODE(clknet_1_0__leaf_net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_B1 (.DIODE(clknet_1_0__leaf_net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A2 (.DIODE(clknet_1_0__leaf_net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_S1 (.DIODE(clknet_1_0__leaf_net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net635_X (.DIODE(clknet_1_0__leaf_net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_S0 (.DIODE(clknet_1_1__leaf_net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A3 (.DIODE(clknet_1_1__leaf_net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(clknet_1_1__leaf_net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A3 (.DIODE(clknet_1_1__leaf_net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net635_X (.DIODE(clknet_1_1__leaf_net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A2 (.DIODE(clknet_1_0__leaf_net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A1 (.DIODE(clknet_1_0__leaf_net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net1003_X (.DIODE(clknet_1_0__leaf_net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A0 (.DIODE(clknet_1_1__leaf_net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A2 (.DIODE(clknet_1_1__leaf_net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A0 (.DIODE(clknet_1_1__leaf_net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net82_X (.DIODE(clknet_1_1__leaf_net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A2 (.DIODE(clknet_1_0__leaf_net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A2 (.DIODE(clknet_1_0__leaf_net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A0 (.DIODE(clknet_1_0__leaf_net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A3 (.DIODE(clknet_1_0__leaf_net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net83_X (.DIODE(clknet_1_0__leaf_net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net979_A (.DIODE(clknet_0_net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net979_A (.DIODE(clknet_0_net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net979_X (.DIODE(clknet_0_net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A1 (.DIODE(clknet_1_0__leaf_net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(clknet_1_0__leaf_net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A2 (.DIODE(clknet_1_0__leaf_net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net979_X (.DIODE(clknet_1_0__leaf_net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A3 (.DIODE(clknet_1_0__leaf_net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A2 (.DIODE(clknet_1_0__leaf_net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_S1 (.DIODE(clknet_1_0__leaf_net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A3 (.DIODE(clknet_1_0__leaf_net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_S0 (.DIODE(clknet_1_0__leaf_net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net704_X (.DIODE(clknet_1_0__leaf_net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_SET_B (.DIODE(clknet_1_1__leaf_net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_S0 (.DIODE(clknet_1_1__leaf_net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S1 (.DIODE(clknet_1_1__leaf_net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S0 (.DIODE(clknet_1_1__leaf_net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net704_X (.DIODE(clknet_1_1__leaf_net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A1 (.DIODE(clknet_1_0__leaf_net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(clknet_1_0__leaf_net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net241_X (.DIODE(clknet_1_0__leaf_net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_S1 (.DIODE(clknet_1_0__leaf_net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S0 (.DIODE(clknet_1_0__leaf_net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_S1 (.DIODE(clknet_1_0__leaf_net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_SET_B (.DIODE(clknet_1_0__leaf_net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A2 (.DIODE(clknet_1_0__leaf_net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S1 (.DIODE(clknet_1_0__leaf_net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_S0 (.DIODE(clknet_1_0__leaf_net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net703_X (.DIODE(clknet_1_0__leaf_net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_S0 (.DIODE(clknet_1_1__leaf_net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_S1 (.DIODE(clknet_1_1__leaf_net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A2 (.DIODE(clknet_1_1__leaf_net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S0 (.DIODE(clknet_1_1__leaf_net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S1 (.DIODE(clknet_1_1__leaf_net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S0 (.DIODE(clknet_1_1__leaf_net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net703_X (.DIODE(clknet_1_1__leaf_net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer3_A (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A3 (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_A (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S0 (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_X (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net1109));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net146),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net1172),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net746),
    .X(net1174));
 sky130_fd_sc_hd__clkbuf_1 clone15 (.A(clknet_0_net255),
    .X(net1175));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
