module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in3,
    in4,
    in5,
    in6,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out3,
    out4,
    out5,
    out6,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in3;
 input in4;
 input in5;
 input in6;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out3;
 output out4;
 output out5;
 output out6;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net631;
 wire net754;
 wire net765;
 wire net770;
 wire net781;
 wire net794;
 wire net811;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_0_net1093;
 wire clknet_1_0__leaf_net1093;
 wire clknet_1_1__leaf_net1093;
 wire clknet_0_net1154;
 wire clknet_1_0__leaf_net1154;
 wire clknet_1_1__leaf_net1154;
 wire clknet_0_net1092;
 wire clknet_1_0__leaf_net1092;
 wire clknet_1_1__leaf_net1092;
 wire clknet_0_net886;
 wire clknet_1_0__leaf_net886;
 wire clknet_1_1__leaf_net886;
 wire clknet_0_net1091;
 wire clknet_1_0__leaf_net1091;
 wire clknet_1_1__leaf_net1091;
 wire clknet_0_net848;
 wire clknet_1_0__leaf_net848;
 wire clknet_1_1__leaf_net848;
 wire clknet_0_net608;
 wire clknet_1_0__leaf_net608;
 wire clknet_1_1__leaf_net608;
 wire clknet_0_net615;
 wire clknet_1_0__leaf_net615;
 wire clknet_1_1__leaf_net615;
 wire clknet_0_net892;
 wire clknet_1_0__leaf_net892;
 wire clknet_1_1__leaf_net892;
 wire clknet_0_net1153;
 wire clknet_1_0__leaf_net1153;
 wire clknet_1_1__leaf_net1153;
 wire clknet_0_net507;
 wire clknet_1_0__leaf_net507;
 wire clknet_1_1__leaf_net507;
 wire clknet_0_net1160;
 wire clknet_1_0__leaf_net1160;
 wire clknet_1_1__leaf_net1160;
 wire clknet_0_net1150;
 wire clknet_1_0__leaf_net1150;
 wire clknet_1_1__leaf_net1150;
 wire clknet_0_net1072;
 wire clknet_1_0__leaf_net1072;
 wire clknet_1_1__leaf_net1072;
 wire clknet_0_net574;
 wire clknet_1_0__leaf_net574;
 wire clknet_1_1__leaf_net574;
 wire clknet_0_net1109;
 wire clknet_1_0__leaf_net1109;
 wire clknet_1_1__leaf_net1109;
 wire clknet_0_net1111;
 wire clknet_1_0__leaf_net1111;
 wire clknet_1_1__leaf_net1111;
 wire clknet_0_net689;
 wire clknet_1_0__leaf_net689;
 wire clknet_1_1__leaf_net689;
 wire clknet_0_net570;
 wire clknet_1_0__leaf_net570;
 wire clknet_1_1__leaf_net570;
 wire clknet_0_net1071;
 wire clknet_1_0__leaf_net1071;
 wire clknet_1_1__leaf_net1071;
 wire clknet_0_net1070;
 wire clknet_1_0__leaf_net1070;
 wire clknet_1_1__leaf_net1070;
 wire clknet_0_net1052;
 wire clknet_1_0__leaf_net1052;
 wire clknet_1_1__leaf_net1052;
 wire clknet_0_net1051;
 wire clknet_1_0__leaf_net1051;
 wire clknet_1_1__leaf_net1051;
 wire clknet_0_net1050;
 wire clknet_1_0__leaf_net1050;
 wire clknet_1_1__leaf_net1050;
 wire clknet_0_net524;
 wire clknet_1_0__leaf_net524;
 wire clknet_1_1__leaf_net524;
 wire clknet_0_net1032;
 wire clknet_1_0__leaf_net1032;
 wire clknet_1_1__leaf_net1032;
 wire clknet_0_net458;
 wire clknet_1_0__leaf_net458;
 wire clknet_1_1__leaf_net458;
 wire clknet_0_net1031;
 wire clknet_1_0__leaf_net1031;
 wire clknet_1_1__leaf_net1031;
 wire clknet_0_net457;
 wire clknet_1_0__leaf_net457;
 wire clknet_1_1__leaf_net457;
 wire clknet_0_net1030;
 wire clknet_1_0__leaf_net1030;
 wire clknet_1_1__leaf_net1030;
 wire clknet_0_net1011;
 wire clknet_1_0__leaf_net1011;
 wire clknet_1_1__leaf_net1011;
 wire clknet_0_net1010;
 wire clknet_1_0__leaf_net1010;
 wire clknet_1_1__leaf_net1010;
 wire clknet_0_net381;
 wire clknet_1_0__leaf_net381;
 wire clknet_1_1__leaf_net381;
 wire clknet_0_net385;
 wire clknet_1_0__leaf_net385;
 wire clknet_1_1__leaf_net385;
 wire clknet_0_net1009;
 wire clknet_1_0__leaf_net1009;
 wire clknet_1_1__leaf_net1009;
 wire clknet_0_net990;
 wire clknet_1_0__leaf_net990;
 wire clknet_1_1__leaf_net990;
 wire clknet_0_net417;
 wire clknet_1_0__leaf_net417;
 wire clknet_1_1__leaf_net417;
 wire clknet_0_net418;
 wire clknet_1_0__leaf_net418;
 wire clknet_1_1__leaf_net418;
 wire clknet_0_net290;
 wire clknet_1_0__leaf_net290;
 wire clknet_1_1__leaf_net290;
 wire clknet_0_net989;
 wire clknet_1_0__leaf_net989;
 wire clknet_1_1__leaf_net989;
 wire clknet_0_net988;
 wire clknet_1_0__leaf_net988;
 wire clknet_1_1__leaf_net988;
 wire clknet_0_net969;
 wire clknet_1_0__leaf_net969;
 wire clknet_1_1__leaf_net969;
 wire clknet_0_net341;
 wire clknet_1_0__leaf_net341;
 wire clknet_1_1__leaf_net341;
 wire clknet_0_net228;
 wire clknet_1_0__leaf_net228;
 wire clknet_1_1__leaf_net228;
 wire clknet_0_net968;
 wire clknet_1_0__leaf_net968;
 wire clknet_1_1__leaf_net968;
 wire clknet_0_net487;
 wire clknet_1_0__leaf_net487;
 wire clknet_1_1__leaf_net487;
 wire clknet_0_net503;
 wire clknet_1_0__leaf_net503;
 wire clknet_1_1__leaf_net503;
 wire clknet_0_net499;
 wire clknet_1_0__leaf_net499;
 wire clknet_1_1__leaf_net499;
 wire clknet_0_net492;
 wire clknet_1_0__leaf_net492;
 wire clknet_1_1__leaf_net492;
 wire clknet_0_net489;
 wire clknet_1_0__leaf_net489;
 wire clknet_1_1__leaf_net489;
 wire clknet_0_net488;
 wire clknet_1_0__leaf_net488;
 wire clknet_1_1__leaf_net488;
 wire clknet_0_net238;
 wire clknet_1_0__leaf_net238;
 wire clknet_1_1__leaf_net238;
 wire clknet_0_net227;
 wire clknet_1_0__leaf_net227;
 wire clknet_1_1__leaf_net227;
 wire clknet_0_net226;
 wire clknet_1_0__leaf_net226;
 wire clknet_1_1__leaf_net226;
 wire clknet_0_net967;
 wire clknet_1_0__leaf_net967;
 wire clknet_1_1__leaf_net967;
 wire clknet_0_net948;
 wire clknet_1_0__leaf_net948;
 wire clknet_1_1__leaf_net948;
 wire clknet_0_net297;
 wire clknet_1_0__leaf_net297;
 wire clknet_1_1__leaf_net297;
 wire clknet_0_net891;
 wire clknet_1_0__leaf_net891;
 wire clknet_1_1__leaf_net891;
 wire clknet_0_net595;
 wire clknet_1_0__leaf_net595;
 wire clknet_1_1__leaf_net595;
 wire clknet_0_net692;
 wire clknet_1_0__leaf_net692;
 wire clknet_1_1__leaf_net692;
 wire clknet_0_net694;
 wire clknet_1_0__leaf_net694;
 wire clknet_1_1__leaf_net694;
 wire clknet_0_net618;
 wire clknet_1_0__leaf_net618;
 wire clknet_1_1__leaf_net618;
 wire clknet_0_net619;
 wire clknet_1_0__leaf_net619;
 wire clknet_1_1__leaf_net619;
 wire clknet_0_net596;
 wire clknet_1_0__leaf_net596;
 wire clknet_1_1__leaf_net596;
 wire clknet_0_net202;
 wire clknet_1_0__leaf_net202;
 wire clknet_1_1__leaf_net202;
 wire clknet_0_net220;
 wire clknet_1_0__leaf_net220;
 wire clknet_1_1__leaf_net220;
 wire clknet_0_net846;
 wire clknet_1_0__leaf_net846;
 wire clknet_1_1__leaf_net846;
 wire clknet_0_net216;
 wire clknet_1_0__leaf_net216;
 wire clknet_1_1__leaf_net216;
 wire clknet_0_net211;
 wire clknet_1_0__leaf_net211;
 wire clknet_1_1__leaf_net211;
 wire clknet_0_net210;
 wire clknet_1_0__leaf_net210;
 wire clknet_1_1__leaf_net210;
 wire clknet_0_net208;
 wire clknet_1_0__leaf_net208;
 wire clknet_1_1__leaf_net208;
 wire clknet_0_net205;
 wire clknet_1_0__leaf_net205;
 wire clknet_1_1__leaf_net205;
 wire clknet_0_net204;
 wire clknet_1_0__leaf_net204;
 wire clknet_1_1__leaf_net204;
 wire clknet_0_net203;
 wire clknet_1_0__leaf_net203;
 wire clknet_1_1__leaf_net203;
 wire clknet_0_net298;
 wire clknet_1_0__leaf_net298;
 wire clknet_1_1__leaf_net298;
 wire clknet_0_net890;
 wire clknet_1_0__leaf_net890;
 wire clknet_1_1__leaf_net890;
 wire clknet_0_net469;
 wire clknet_1_0__leaf_net469;
 wire clknet_1_1__leaf_net469;
 wire clknet_0_net483;
 wire clknet_1_0__leaf_net483;
 wire clknet_1_1__leaf_net483;
 wire clknet_0_net479;
 wire clknet_1_0__leaf_net479;
 wire clknet_1_1__leaf_net479;
 wire clknet_0_net482;
 wire clknet_1_0__leaf_net482;
 wire clknet_1_1__leaf_net482;
 wire clknet_0_net465;
 wire clknet_1_0__leaf_net465;
 wire clknet_1_1__leaf_net465;
 wire clknet_0_net947;
 wire clknet_1_0__leaf_net947;
 wire clknet_1_1__leaf_net947;
 wire clknet_0_net200;
 wire clknet_1_0__leaf_net200;
 wire clknet_1_1__leaf_net200;
 wire clknet_0_net318;
 wire clknet_1_0__leaf_net318;
 wire clknet_1_1__leaf_net318;
 wire clknet_0_net180;
 wire clknet_1_0__leaf_net180;
 wire clknet_1_1__leaf_net180;
 wire clknet_0_net195;
 wire clknet_1_0__leaf_net195;
 wire clknet_1_1__leaf_net195;
 wire clknet_0_net185;
 wire clknet_1_0__leaf_net185;
 wire clknet_1_1__leaf_net185;
 wire clknet_0_net181;
 wire clknet_1_0__leaf_net181;
 wire clknet_1_1__leaf_net181;
 wire clknet_0_net179;
 wire clknet_1_0__leaf_net179;
 wire clknet_1_1__leaf_net179;
 wire clknet_0_net946;
 wire clknet_1_0__leaf_net946;
 wire clknet_1_1__leaf_net946;
 wire clknet_0_net927;
 wire clknet_1_0__leaf_net927;
 wire clknet_1_1__leaf_net927;
 wire clknet_0_net248;
 wire clknet_1_0__leaf_net248;
 wire clknet_1_1__leaf_net248;
 wire clknet_0_net260;
 wire clknet_1_0__leaf_net260;
 wire clknet_1_1__leaf_net260;
 wire clknet_0_net252;
 wire clknet_1_0__leaf_net252;
 wire clknet_1_1__leaf_net252;
 wire clknet_0_net249;
 wire clknet_1_0__leaf_net249;
 wire clknet_1_1__leaf_net249;
 wire clknet_0_net247;
 wire clknet_1_0__leaf_net247;
 wire clknet_1_1__leaf_net247;
 wire clknet_0_net127;
 wire clknet_1_0__leaf_net127;
 wire clknet_1_1__leaf_net127;
 wire clknet_0_net926;
 wire clknet_1_0__leaf_net926;
 wire clknet_1_1__leaf_net926;
 wire clknet_0_net925;
 wire clknet_1_0__leaf_net925;
 wire clknet_1_1__leaf_net925;
 wire clknet_0_net105;
 wire clknet_1_0__leaf_net105;
 wire clknet_1_1__leaf_net105;
 wire clknet_0_net906;
 wire clknet_1_0__leaf_net906;
 wire clknet_1_1__leaf_net906;
 wire clknet_0_net37;
 wire clknet_1_0__leaf_net37;
 wire clknet_1_1__leaf_net37;
 wire clknet_0_net35;
 wire clknet_1_0__leaf_net35;
 wire clknet_1_1__leaf_net35;
 wire clknet_0_net905;
 wire clknet_1_0__leaf_net905;
 wire clknet_1_1__leaf_net905;
 wire clknet_0_net157;
 wire clknet_1_0__leaf_net157;
 wire clknet_1_1__leaf_net157;
 wire clknet_0_net155;
 wire clknet_1_0__leaf_net155;
 wire clknet_1_1__leaf_net155;
 wire clknet_0_net171;
 wire clknet_1_0__leaf_net171;
 wire clknet_1_1__leaf_net171;
 wire clknet_0_net159;
 wire clknet_1_0__leaf_net159;
 wire clknet_1_1__leaf_net159;
 wire clknet_0_net156;
 wire clknet_1_0__leaf_net156;
 wire clknet_1_1__leaf_net156;
 wire clknet_0_net904;
 wire clknet_1_0__leaf_net904;
 wire clknet_1_1__leaf_net904;
 wire clknet_0_net1128;
 wire clknet_1_0__leaf_net1128;
 wire clknet_1_1__leaf_net1128;
 wire clknet_0_net533;
 wire clknet_1_0__leaf_net533;
 wire clknet_1_1__leaf_net533;
 wire clknet_0_net548;
 wire clknet_1_0__leaf_net548;
 wire clknet_1_1__leaf_net548;
 wire clknet_0_net667;
 wire clknet_1_0__leaf_net667;
 wire clknet_1_1__leaf_net667;
 wire clknet_0_net681;
 wire clknet_1_0__leaf_net681;
 wire clknet_1_1__leaf_net681;
 wire clknet_0_net1110;
 wire clknet_1_0__leaf_net1110;
 wire clknet_1_1__leaf_net1110;
 wire clknet_0_net668;
 wire clknet_1_0__leaf_net668;
 wire clknet_1_1__leaf_net668;
 wire clknet_0_net641;
 wire clknet_1_0__leaf_net641;
 wire clknet_1_1__leaf_net641;
 wire clknet_0_net642;
 wire clknet_1_0__leaf_net642;
 wire clknet_1_1__leaf_net642;
 wire clknet_0_net553;
 wire clknet_1_0__leaf_net553;
 wire clknet_1_1__leaf_net553;
 wire clknet_0_net554;
 wire clknet_1_0__leaf_net554;
 wire clknet_1_1__leaf_net554;
 wire clknet_0_net549;
 wire clknet_1_0__leaf_net549;
 wire clknet_1_1__leaf_net549;
 wire clknet_0_net550;
 wire clknet_1_0__leaf_net550;
 wire clknet_1_1__leaf_net550;
 wire clknet_0_net535;
 wire clknet_1_0__leaf_net535;
 wire clknet_1_1__leaf_net535;
 wire clknet_0_net539;
 wire clknet_1_0__leaf_net539;
 wire clknet_1_1__leaf_net539;
 wire clknet_0_net278;
 wire clknet_1_0__leaf_net278;
 wire clknet_1_1__leaf_net278;
 wire clknet_0_net855;
 wire clknet_1_0__leaf_net855;
 wire clknet_1_1__leaf_net855;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;

 sky130_fd_sc_hd__mux4_1 c100 (.A0(net77),
    .A1(net73),
    .A2(net64),
    .A3(net69),
    .S0(net917),
    .S1(net919),
    .X(net79));
 sky130_fd_sc_hd__mux4_1 c101 (.A0(net70),
    .A1(net65),
    .A2(net69),
    .A3(net917),
    .S0(net919),
    .S1(net920),
    .X(net80));
 sky130_fd_sc_hd__mux4_1 c102 (.A0(net80),
    .A1(net77),
    .A2(net65),
    .A3(net917),
    .S0(net918),
    .S1(net920),
    .X(net81));
 sky130_fd_sc_hd__mux4_1 c103 (.A0(net71),
    .A1(net80),
    .A2(net73),
    .A3(net884),
    .S0(net919),
    .S1(net921),
    .X(net82));
 sky130_fd_sc_hd__mux4_1 c104 (.A0(net80),
    .A1(net76),
    .A2(net884),
    .A3(net917),
    .S0(net918),
    .S1(net921),
    .X(net83));
 sky130_fd_sc_hd__buf_1 c105 (.X(net768));
 sky130_fd_sc_hd__and2_0 c106 (.A(net59),
    .B(net84),
    .X(net85));
 sky130_fd_sc_hd__and2_1 c107 (.A(net72),
    .B(net84),
    .X(net86));
 sky130_fd_sc_hd__and2_1 c108 (.A(net84),
    .B(net1170),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 c109 (.A(net767),
    .X(net88));
 sky130_fd_sc_hd__and2_1 c110 (.A(net88),
    .B(net84),
    .X(net89));
 sky130_fd_sc_hd__sdfbbn_1 c111 (.CLK_N(clknet_leaf_46_clk),
    .D(net1179),
    .RESET_B(net85),
    .SCD(net84),
    .SCE(net88),
    .SET_B(net87),
    .Q(net91),
    .Q_N(net90));
 sky130_fd_sc_hd__mux4_1 c112 (.A0(net91),
    .A1(net60),
    .A2(net1179),
    .A3(net84),
    .S0(net86),
    .S1(net1170),
    .X(net92));
 sky130_fd_sc_hd__or4bb_2 c113 (.A(net1179),
    .B(net91),
    .C_N(net84),
    .D_N(net922),
    .X(net93));
 sky130_fd_sc_hd__a2111o_1 c114 (.A1(net93),
    .A2(net1179),
    .B1(net84),
    .C1(net90),
    .D1(net922),
    .X(net94));
 sky130_fd_sc_hd__sdfbbp_1 c115 (.CLK(clknet_leaf_45_clk),
    .D(net85),
    .RESET_B(net1179),
    .SCD(net84),
    .SCE(net91),
    .SET_B(net1243),
    .Q(net96),
    .Q_N(net95));
 sky130_fd_sc_hd__a2111o_1 c116 (.A1(net95),
    .A2(net84),
    .B1(net1179),
    .C1(net90),
    .D1(net922),
    .X(net97));
 sky130_fd_sc_hd__a2111o_1 c117 (.A1(net96),
    .A2(net93),
    .B1(net97),
    .C1(net1179),
    .D1(net84),
    .X(net98));
 sky130_fd_sc_hd__a2111o_1 c118 (.A1(net97),
    .A2(net1179),
    .B1(net98),
    .C1(net84),
    .D1(net95),
    .X(net99));
 sky130_fd_sc_hd__mux4_2 c119 (.A0(net84),
    .A1(net96),
    .A2(net93),
    .A3(net97),
    .S0(net89),
    .S1(net922),
    .X(net100));
 sky130_fd_sc_hd__mux4_1 c120 (.A0(net94),
    .A1(net98),
    .A2(net100),
    .A3(net97),
    .S0(net95),
    .S1(net922),
    .X(net101));
 sky130_fd_sc_hd__mux4_1 c121 (.A0(net100),
    .A1(net96),
    .A2(net98),
    .A3(net97),
    .S0(net1179),
    .S1(net923),
    .X(net102));
 sky130_fd_sc_hd__mux4_1 c122 (.A0(net97),
    .A1(net85),
    .A2(net100),
    .A3(net841),
    .S0(net923),
    .S1(net924),
    .X(net103));
 sky130_fd_sc_hd__mux4_1 c123 (.A0(net98),
    .A1(net100),
    .A2(net1179),
    .A3(net923),
    .S0(net924),
    .S1(clknet_1_0__leaf_net925),
    .X(net104));
 sky130_fd_sc_hd__mux4_1 c124 (.A0(net59),
    .A1(net841),
    .A2(net884),
    .A3(net923),
    .S0(net924),
    .S1(clknet_1_0__leaf_net925),
    .X(net105));
 sky130_fd_sc_hd__mux4_1 c125 (.A0(clknet_1_0__leaf_net105),
    .A1(net100),
    .A2(net841),
    .A3(net923),
    .S0(net924),
    .S1(clknet_1_1__leaf_net925),
    .X(net106));
 sky130_fd_sc_hd__and2_0 c126 (.A(net1145),
    .B(net1146),
    .X(net107));
 sky130_fd_sc_hd__and2_1 c127 (.A(net1207),
    .B(net765),
    .X(net108));
 sky130_fd_sc_hd__and2_1 c128 (.A(net108),
    .B(net811),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 c129 (.A(net774),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 c130 (.A(net797),
    .X(net111));
 sky130_fd_sc_hd__or4bb_1 c131 (.A(net108),
    .B(net1132),
    .C_N(net109),
    .D_N(net1207),
    .X(net112));
 sky130_fd_sc_hd__and3_1 c132 (.A(net1207),
    .B(net1141),
    .C(net111),
    .X(net113));
 sky130_fd_sc_hd__and3_1 c133 (.A(net113),
    .B(net1208),
    .C(net826),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 c134 (.A(net774),
    .X(net115));
 sky130_fd_sc_hd__sdfbbn_1 c135 (.CLK_N(clknet_leaf_2_clk),
    .D(net111),
    .RESET_B(net113),
    .SCD(net109),
    .SCE(net1207),
    .SET_B(net114),
    .Q(net117),
    .Q_N(net116));
 sky130_fd_sc_hd__buf_1 c136 (.A(net796),
    .X(net118));
 sky130_fd_sc_hd__or4bb_1 c137 (.A(net114),
    .B(net1146),
    .C_N(net111),
    .D_N(net1207),
    .X(net119));
 sky130_fd_sc_hd__and3_1 c138 (.A(net1207),
    .B(net111),
    .C(clknet_1_1__leaf_net855),
    .X(net120));
 sky130_fd_sc_hd__a2111o_1 c139 (.A1(net118),
    .A2(net1207),
    .B1(net113),
    .C1(net111),
    .D1(net116),
    .X(net121));
 sky130_fd_sc_hd__sdfrbp_1 c140 (.CLK(clknet_leaf_10_clk),
    .D(net108),
    .RESET_B(net117),
    .SCD(net121),
    .SCE(net1207),
    .Q(net123),
    .Q_N(net122));
 sky130_fd_sc_hd__mux4_1 c141 (.A0(net111),
    .A1(net123),
    .A2(net121),
    .A3(net1208),
    .S0(net113),
    .S1(clknet_1_1__leaf_net855),
    .X(net124));
 sky130_fd_sc_hd__mux4_1 c142 (.A0(net110),
    .A1(net114),
    .A2(net121),
    .A3(net1207),
    .S0(net118),
    .S1(clknet_1_0__leaf_net927),
    .X(net125));
 sky130_fd_sc_hd__mux4_1 c143 (.A0(net770),
    .A1(net1143),
    .A2(net121),
    .A3(net122),
    .S0(net826),
    .S1(clknet_1_0__leaf_net927),
    .X(net126));
 sky130_fd_sc_hd__mux4_1 c144 (.A0(net115),
    .A1(net123),
    .A2(net1208),
    .A3(net111),
    .S0(clknet_1_0__leaf_net927),
    .S1(net929),
    .X(net127));
 sky130_fd_sc_hd__mux4_1 c145 (.A0(clknet_1_0__leaf_net127),
    .A1(net121),
    .A2(net111),
    .A3(net1208),
    .S0(clknet_1_1__leaf_net927),
    .S1(net929),
    .X(net128));
 sky130_fd_sc_hd__mux4_1 c146 (.A0(net120),
    .A1(net121),
    .A2(clknet_1_1__leaf_net127),
    .A3(clknet_1_0__leaf_net927),
    .S0(net928),
    .S1(net931),
    .X(net129));
 sky130_fd_sc_hd__and2_2 c147 (.A(net1203),
    .B(net930),
    .X(net130));
 sky130_fd_sc_hd__and2_1 c148 (.A(net130),
    .B(net1235),
    .X(net131));
 sky130_fd_sc_hd__and2_0 c149 (.A(net131),
    .B(net130),
    .X(net132));
 sky130_fd_sc_hd__and2_2 c150 (.A(net131),
    .B(net130),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 c151 (.A(net832),
    .X(net134));
 sky130_fd_sc_hd__sdfrbp_1 c152 (.CLK(clknet_leaf_9_clk),
    .D(net130),
    .RESET_B(net131),
    .SCD(net133),
    .SCE(net1204),
    .Q(net136),
    .Q_N(net135));
 sky130_fd_sc_hd__sdfbbn_1 c153 (.CLK_N(clknet_leaf_9_clk),
    .D(net134),
    .RESET_B(net132),
    .SCD(net133),
    .SCE(net130),
    .SET_B(net1204),
    .Q(net138),
    .Q_N(net137));
 sky130_fd_sc_hd__clkbuf_2 c154 (.A(net832),
    .X(net139));
 sky130_fd_sc_hd__sdfbbp_1 c155 (.CLK(clknet_leaf_9_clk),
    .D(net1245),
    .RESET_B(net137),
    .SCD(net139),
    .SCE(net133),
    .SET_B(net130),
    .Q(net141),
    .Q_N(net140));
 sky130_fd_sc_hd__sdfbbn_1 c156 (.CLK_N(clknet_leaf_2_clk),
    .D(net1253),
    .RESET_B(net133),
    .SCD(net141),
    .SCE(net139),
    .SET_B(net131),
    .Q(net143),
    .Q_N(net142));
 sky130_fd_sc_hd__mux4_1 c157 (.A0(net143),
    .A1(net141),
    .A2(net130),
    .A3(net133),
    .S0(net139),
    .S1(net1203),
    .X(net144));
 sky130_fd_sc_hd__mux4_1 c158 (.A0(net133),
    .A1(net141),
    .A2(net143),
    .A3(net139),
    .S0(net130),
    .S1(net934),
    .X(net145));
 sky130_fd_sc_hd__mux4_1 c159 (.A0(net131),
    .A1(net132),
    .A2(net133),
    .A3(net139),
    .S0(net933),
    .S1(net935),
    .X(net146));
 sky130_fd_sc_hd__mux4_1 c160 (.A0(net141),
    .A1(net143),
    .A2(net139),
    .A3(net130),
    .S0(net935),
    .S1(net936),
    .X(net147));
 sky130_fd_sc_hd__mux4_2 c161 (.A0(net136),
    .A1(net147),
    .A2(net140),
    .A3(net142),
    .S0(net935),
    .S1(net936),
    .X(net148));
 sky130_fd_sc_hd__mux4_1 c162 (.A0(net147),
    .A1(net138),
    .A2(net148),
    .A3(net142),
    .S0(net140),
    .S1(net1274),
    .X(net149));
 sky130_fd_sc_hd__mux4_1 c163 (.A0(net147),
    .A1(net148),
    .A2(net140),
    .A3(net1204),
    .S0(net934),
    .S1(net1275),
    .X(net150));
 sky130_fd_sc_hd__mux4_1 c164 (.A0(net135),
    .A1(net134),
    .A2(net147),
    .A3(net139),
    .S0(net148),
    .S1(net938),
    .X(net151));
 sky130_fd_sc_hd__mux4_1 c165 (.A0(net148),
    .A1(net139),
    .A2(net936),
    .A3(net937),
    .S0(net938),
    .S1(net940),
    .X(net152));
 sky130_fd_sc_hd__mux4_1 c166 (.A0(net134),
    .A1(net1140),
    .A2(net139),
    .A3(net833),
    .S0(net938),
    .S1(net939),
    .X(net153));
 sky130_fd_sc_hd__mux4_1 c167 (.A0(net139),
    .A1(net142),
    .A2(net833),
    .A3(net935),
    .S0(net938),
    .S1(net940),
    .X(net154));
 sky130_fd_sc_hd__and2_0 c168 (.A(net865),
    .B(clknet_1_0__leaf_net905),
    .X(net155));
 sky130_fd_sc_hd__and2_0 c169 (.A(clknet_1_1__leaf_net155),
    .B(net1203),
    .X(net156));
 sky130_fd_sc_hd__and3_1 c170 (.A(clknet_1_1__leaf_net156),
    .B(clknet_1_0__leaf_net905),
    .C(net909),
    .X(net157));
 sky130_fd_sc_hd__buf_1 c171 (.A(net785),
    .X(net158));
 sky130_fd_sc_hd__and3_1 c172 (.A(net158),
    .B(clknet_1_1__leaf_net155),
    .C(clknet_1_1__leaf_net156),
    .X(net159));
 sky130_fd_sc_hd__sdfbbn_2 c173 (.CLK_N(clknet_leaf_3_clk),
    .D(clknet_1_0__leaf_net159),
    .RESET_B(net1217),
    .SCD(clknet_1_1__leaf_net156),
    .SCE(clknet_1_1__leaf_net155),
    .SET_B(clknet_1_1__leaf_net905),
    .Q(net161),
    .Q_N(net160));
 sky130_fd_sc_hd__mux4_1 c174 (.A0(net161),
    .A1(net154),
    .A2(clknet_1_0__leaf_net159),
    .A3(clknet_1_1__leaf_net155),
    .S0(clknet_1_1__leaf_net156),
    .S1(net932),
    .X(net162));
 sky130_fd_sc_hd__sdfbbp_1 c175 (.CLK(clknet_leaf_3_clk),
    .D(clknet_1_0__leaf_net155),
    .RESET_B(net1217),
    .SCD(clknet_1_0__leaf_net159),
    .SCE(net160),
    .SET_B(net910),
    .Q(net164),
    .Q_N(net163));
 sky130_fd_sc_hd__sdfbbn_1 c176 (.CLK_N(clknet_leaf_3_clk),
    .D(clknet_1_1__leaf_net156),
    .RESET_B(net164),
    .SCD(clknet_1_0__leaf_net159),
    .SCE(net161),
    .SET_B(clknet_1_0__leaf_net157),
    .Q(net166),
    .Q_N(net165));
 sky130_fd_sc_hd__mux4_1 c177 (.A0(net161),
    .A1(net163),
    .A2(clknet_1_0__leaf_net159),
    .A3(clknet_1_0__leaf_net155),
    .S0(net908),
    .S1(net931),
    .X(net167));
 sky130_fd_sc_hd__mux4_1 c178 (.A0(net165),
    .A1(net164),
    .A2(net160),
    .A3(clknet_1_1__leaf_net159),
    .S0(net813),
    .S1(net941),
    .X(net168));
 sky130_fd_sc_hd__mux4_1 c179 (.A0(net166),
    .A1(net161),
    .A2(net163),
    .A3(clknet_1_1__leaf_net159),
    .S0(clknet_1_0__leaf_net156),
    .S1(net943),
    .X(net169));
 sky130_fd_sc_hd__mux4_1 c180 (.A0(clknet_1_1__leaf_net159),
    .A1(net164),
    .A2(clknet_1_0__leaf_net156),
    .A3(net160),
    .S0(net941),
    .S1(net944),
    .X(net170));
 sky130_fd_sc_hd__mux4_1 c181 (.A0(clknet_1_0__leaf_net155),
    .A1(clknet_1_1__leaf_net156),
    .A2(net163),
    .A3(net160),
    .S0(net942),
    .S1(net943),
    .X(net171));
 sky130_fd_sc_hd__mux4_1 c182 (.A0(net164),
    .A1(clknet_1_1__leaf_net159),
    .A2(clknet_1_1__leaf_net171),
    .A3(net160),
    .S0(clknet_1_0__leaf_net156),
    .S1(net945),
    .X(net172));
 sky130_fd_sc_hd__mux4_1 c183 (.A0(net161),
    .A1(clknet_1_0__leaf_net171),
    .A2(clknet_1_1__leaf_net159),
    .A3(net943),
    .S0(net944),
    .S1(clknet_1_1__leaf_net946),
    .X(net173));
 sky130_fd_sc_hd__mux4_1 c184 (.A0(clknet_1_0__leaf_net156),
    .A1(net161),
    .A2(clknet_1_1__leaf_net171),
    .A3(net944),
    .S0(clknet_1_0__leaf_net946),
    .S1(clknet_1_1__leaf_net947),
    .X(net174));
 sky130_fd_sc_hd__mux4_1 c185 (.A0(clknet_1_0__leaf_net156),
    .A1(clknet_1_1__leaf_net159),
    .A2(net161),
    .A3(clknet_1_1__leaf_net171),
    .S0(net942),
    .S1(clknet_1_1__leaf_net946),
    .X(net175));
 sky130_fd_sc_hd__mux4_1 c186 (.A0(clknet_1_1__leaf_net171),
    .A1(net943),
    .A2(net944),
    .A3(clknet_1_0__leaf_net946),
    .S0(clknet_1_1__leaf_net947),
    .S1(clknet_1_0__leaf_net948),
    .X(net176));
 sky130_fd_sc_hd__mux4_1 c187 (.A0(net158),
    .A1(clknet_1_1__leaf_net159),
    .A2(clknet_1_1__leaf_net171),
    .A3(net160),
    .S0(clknet_1_0__leaf_net890),
    .S1(clknet_1_0__leaf_net948),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 c188 (.A0(net153),
    .A1(clknet_1_1__leaf_net171),
    .A2(net813),
    .A3(clknet_1_0__leaf_net890),
    .S0(net945),
    .S1(net949),
    .X(net178));
 sky130_fd_sc_hd__and2_0 c189 (.A(net880),
    .B(clknet_1_1__leaf_net947),
    .X(net179));
 sky130_fd_sc_hd__and2_0 c190 (.A(clknet_1_0__leaf_net179),
    .B(clknet_1_0__leaf_net947),
    .X(net180));
 sky130_fd_sc_hd__and2_0 c191 (.A(clknet_1_0__leaf_net180),
    .B(clknet_1_0__leaf_net179),
    .X(net181));
 sky130_fd_sc_hd__sdfrtn_1 c192 (.CLK_N(clknet_leaf_3_clk),
    .D(clknet_1_0__leaf_net181),
    .RESET_B(clknet_1_0__leaf_net179),
    .SCD(net908),
    .SCE(clknet_1_0__leaf_net947),
    .Q(net182));
 sky130_fd_sc_hd__sdfbbn_1 c193 (.CLK_N(clknet_leaf_0_clk),
    .D(clknet_1_0__leaf_net171),
    .RESET_B(net182),
    .SCD(clknet_1_0__leaf_net180),
    .SCE(clknet_1_0__leaf_net179),
    .SET_B(clknet_1_0__leaf_net947),
    .Q(net184),
    .Q_N(net183));
 sky130_fd_sc_hd__a2111o_1 c194 (.A1(net184),
    .A2(clknet_1_0__leaf_net179),
    .B1(net182),
    .C1(clknet_1_0__leaf_net180),
    .D1(net842),
    .X(net185));
 sky130_fd_sc_hd__mux4_1 c195 (.A0(clknet_1_0__leaf_net181),
    .A1(clknet_1_0__leaf_net171),
    .A2(clknet_1_0__leaf_net185),
    .A3(net183),
    .S0(clknet_1_0__leaf_net180),
    .S1(clknet_1_0__leaf_net179),
    .X(net186));
 sky130_fd_sc_hd__mux4_1 c196 (.A0(clknet_1_0__leaf_net180),
    .A1(net182),
    .A2(clknet_1_0__leaf_net185),
    .A3(clknet_1_0__leaf_net179),
    .S0(net183),
    .S1(net952),
    .X(net187));
 sky130_fd_sc_hd__mux4_1 c197 (.A0(clknet_1_0__leaf_net185),
    .A1(clknet_1_0__leaf_net171),
    .A2(net844),
    .A3(net865),
    .S0(clknet_1_0__leaf_net947),
    .S1(net952),
    .X(net188));
 sky130_fd_sc_hd__mux4_1 c198 (.A0(clknet_1_0__leaf_net185),
    .A1(net183),
    .A2(net182),
    .A3(clknet_1_1__leaf_net179),
    .S1(net953),
    .X(net189));
 sky130_fd_sc_hd__mux4_1 c199 (.A0(net184),
    .A1(clknet_1_1__leaf_net180),
    .A2(clknet_1_1__leaf_net185),
    .A3(clknet_1_1__leaf_net179),
    .S0(net952),
    .S1(net954),
    .X(net190));
 sky130_fd_sc_hd__mux4_1 c200 (.A0(clknet_1_0__leaf_net179),
    .A1(clknet_1_0__leaf_net185),
    .A2(net843),
    .A3(net907),
    .S0(net951),
    .S1(net954),
    .X(net191));
 sky130_fd_sc_hd__mux4_1 c201 (.A0(clknet_1_0__leaf_net185),
    .A1(clknet_1_1__leaf_net180),
    .A2(clknet_1_0__leaf_net171),
    .A3(clknet_1_1__leaf_net179),
    .S0(net953),
    .S1(net956),
    .X(net192));
 sky130_fd_sc_hd__mux4_1 c202 (.A0(clknet_1_1__leaf_net180),
    .A1(clknet_1_1__leaf_net185),
    .A2(net951),
    .A3(net954),
    .S0(net955),
    .S1(net957),
    .X(net193));
 sky130_fd_sc_hd__mux4_1 c203 (.A0(net182),
    .A1(clknet_1_1__leaf_net185),
    .A2(net952),
    .A3(net953),
    .S0(net957),
    .S1(net958),
    .X(net194));
 sky130_fd_sc_hd__mux4_1 c204 (.A0(clknet_1_1__leaf_net180),
    .A1(clknet_1_1__leaf_net179),
    .A2(net844),
    .A3(net951),
    .S0(net956),
    .S1(net959),
    .X(net195));
 sky130_fd_sc_hd__mux4_1 c205 (.A0(clknet_1_0__leaf_net181),
    .A1(clknet_1_1__leaf_net179),
    .A2(net954),
    .A3(net955),
    .S0(net957),
    .S1(net958),
    .X(net196));
 sky130_fd_sc_hd__mux4_1 c206 (.A0(clknet_1_0__leaf_net195),
    .A1(net183),
    .A2(net956),
    .A3(net958),
    .S0(net959),
    .S1(net960),
    .X(net197));
 sky130_fd_sc_hd__mux4_1 c207 (.A0(clknet_1_1__leaf_net195),
    .A1(clknet_1_1__leaf_net185),
    .A2(net182),
    .A3(net958),
    .S0(net961),
    .S1(net962),
    .X(net198));
 sky130_fd_sc_hd__mux4_1 c208 (.A0(net953),
    .A1(net955),
    .A2(net959),
    .A3(net961),
    .S0(net963),
    .S1(net964),
    .X(net199));
 sky130_fd_sc_hd__mux4_1 c209 (.A0(net199),
    .A1(clknet_1_1__leaf_net947),
    .A2(net958),
    .A3(net960),
    .S0(net963),
    .S1(net964),
    .X(net200));
 sky130_fd_sc_hd__and2_1 c210 (.A(net1171),
    .B(net964),
    .X(net201));
 sky130_fd_sc_hd__and2_0 c211 (.A(net62),
    .B(clknet_1_0__leaf_net891),
    .X(net202));
 sky130_fd_sc_hd__and2_0 c212 (.A(net1167),
    .B(clknet_1_1__leaf_net202),
    .X(net203));
 sky130_fd_sc_hd__and3_1 c213 (.A(net184),
    .B(clknet_1_1__leaf_net202),
    .C(net1167),
    .X(net204));
 sky130_fd_sc_hd__a2111o_1 c214 (.A1(net1171),
    .A2(clknet_1_1__leaf_net202),
    .B1(net1167),
    .C1(clknet_1_0__leaf_net204),
    .D1(net964),
    .X(net205));
 sky130_fd_sc_hd__buf_1 c215 (.A(net894),
    .X(net206));
 sky130_fd_sc_hd__sdfrtp_1 c216 (.CLK(clknet_leaf_43_clk),
    .D(clknet_1_1__leaf_net204),
    .RESET_B(clknet_1_1__leaf_net202),
    .SCD(clknet_1_1__leaf_net181),
    .SCE(clknet_1_0__leaf_net205),
    .Q(net207));
 sky130_fd_sc_hd__and3_1 c217 (.A(net206),
    .B(net1167),
    .C(clknet_1_0__leaf_net202),
    .X(net208));
 sky130_fd_sc_hd__or4bb_1 c218 (.A(clknet_1_1__leaf_net208),
    .B(net1167),
    .C_N(clknet_1_1__leaf_net202),
    .D_N(clknet_1_0__leaf_net205),
    .X(net209));
 sky130_fd_sc_hd__or4bb_1 c219 (.A(net207),
    .B(clknet_1_0__leaf_net202),
    .C_N(clknet_1_0__leaf_net208),
    .D_N(net1167),
    .X(net210));
 sky130_fd_sc_hd__a2111o_1 c220 (.A1(net207),
    .A2(clknet_1_0__leaf_net208),
    .B1(clknet_1_0__leaf_net202),
    .C1(net1168),
    .D1(net206),
    .X(net211));
 sky130_fd_sc_hd__sdfbbp_1 c221 (.CLK(clknet_leaf_44_clk),
    .D(clknet_1_1__leaf_net210),
    .RESET_B(net207),
    .SCD(clknet_1_0__leaf_net208),
    .SCE(net1167),
    .SET_B(clknet_1_0__leaf_net202),
    .Q(net213),
    .Q_N(net212));
 sky130_fd_sc_hd__sdfbbn_2 c222 (.CLK_N(clknet_leaf_45_clk),
    .D(net213),
    .RESET_B(clknet_1_0__leaf_net208),
    .SCD(clknet_1_0__leaf_net210),
    .SCE(clknet_1_0__leaf_net202),
    .SET_B(net1167),
    .Q(net215),
    .Q_N(net214));
 sky130_fd_sc_hd__mux4_1 c223 (.A0(clknet_1_1__leaf_net202),
    .A1(clknet_1_0__leaf_net208),
    .A2(net214),
    .A3(net1167),
    .S0(net207),
    .S1(clknet_1_1__leaf_net846),
    .X(net216));
 sky130_fd_sc_hd__mux4_1 c224 (.A0(clknet_1_0__leaf_net203),
    .A1(net1168),
    .A2(net215),
    .A3(clknet_1_1__leaf_net208),
    .S0(clknet_1_1__leaf_net202),
    .S1(clknet_1_1__leaf_net216),
    .X(net217));
 sky130_fd_sc_hd__mux4_1 c225 (.A0(clknet_1_0__leaf_net211),
    .A1(net215),
    .A2(clknet_1_1__leaf_net208),
    .A3(clknet_1_0__leaf_net202),
    .S0(net1171),
    .S1(clknet_1_0__leaf_net846),
    .X(net218));
 sky130_fd_sc_hd__mux4_1 c226 (.A0(clknet_1_1__leaf_net211),
    .A1(net215),
    .A2(clknet_1_1__leaf_net208),
    .A3(clknet_1_0__leaf_net202),
    .S0(net1168),
    .S1(clknet_1_0__leaf_net846),
    .X(net219));
 sky130_fd_sc_hd__mux4_1 c227 (.A0(clknet_1_0__leaf_net208),
    .A1(net1167),
    .A2(net214),
    .A3(net212),
    .S0(clknet_1_0__leaf_net202),
    .S1(net965),
    .X(net220));
 sky130_fd_sc_hd__mux4_1 c228 (.A0(clknet_1_0__leaf_net220),
    .A1(net213),
    .A2(net184),
    .A3(net1171),
    .S0(clknet_1_1__leaf_net846),
    .S1(net966),
    .X(net221));
 sky130_fd_sc_hd__mux4_1 c229 (.A0(clknet_1_1__leaf_net205),
    .A1(clknet_1_0__leaf_net220),
    .A2(net214),
    .A3(clknet_1_1__leaf_net208),
    .S0(net1168),
    .S1(clknet_1_1__leaf_net967),
    .X(net222));
 sky130_fd_sc_hd__mux4_1 c230 (.A0(clknet_1_0__leaf_net216),
    .A1(clknet_1_1__leaf_net220),
    .A2(net965),
    .A3(net966),
    .S0(clknet_1_0__leaf_net967),
    .S1(clknet_1_1__leaf_net968),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_2 c231 (.X(net224));
 sky130_fd_sc_hd__buf_2 c232 (.A(net780),
    .X(net225));
 sky130_fd_sc_hd__a2111o_1 c233 (.A1(net215),
    .A2(net225),
    .B1(net224),
    .C1(clknet_1_1__leaf_net926),
    .D1(clknet_1_0__leaf_net968),
    .X(net226));
 sky130_fd_sc_hd__or4bb_1 c234 (.A(clknet_1_1__leaf_net226),
    .B(net225),
    .C_N(net224),
    .D_N(clknet_1_0__leaf_net968),
    .X(net227));
 sky130_fd_sc_hd__and3_1 c235 (.A(clknet_1_1__leaf_net227),
    .B(net225),
    .C(clknet_1_0__leaf_net969),
    .X(net228));
 sky130_fd_sc_hd__sdfbbn_1 c236 (.CLK_N(clknet_leaf_39_clk),
    .D(clknet_1_0__leaf_net228),
    .RESET_B(net1218),
    .SCD(clknet_1_0__leaf_net105),
    .SCE(clknet_1_0__leaf_net227),
    .SET_B(clknet_1_0__leaf_net926),
    .Q(net230),
    .Q_N(net229));
 sky130_fd_sc_hd__a2111o_1 c237 (.A1(net224),
    .A2(clknet_1_1__leaf_net227),
    .B1(net230),
    .C1(clknet_1_0__leaf_net228),
    .D1(net225),
    .X(net231));
 sky130_fd_sc_hd__a2111o_1 c238 (.A1(net1216),
    .A2(clknet_1_1__leaf_net228),
    .B1(clknet_1_0__leaf_net105),
    .C1(clknet_1_1__leaf_net227),
    .D1(clknet_1_0__leaf_net969),
    .X(net232));
 sky130_fd_sc_hd__sdfbbp_1 c239 (.CLK(clknet_leaf_39_clk),
    .D(clknet_1_0__leaf_net226),
    .RESET_B(clknet_1_0__leaf_net227),
    .SCD(net229),
    .SCE(clknet_1_0__leaf_net228),
    .SET_B(net1216),
    .Q(net234),
    .Q_N(net233));
 sky130_fd_sc_hd__a2111o_1 c240 (.A1(net230),
    .A2(net234),
    .B1(clknet_1_0__leaf_net228),
    .C1(clknet_1_0__leaf_net226),
    .D1(clknet_1_0__leaf_net227),
    .X(net235));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(net230),
    .A1(net234),
    .A2(clknet_1_0__leaf_net227),
    .A3(net225),
    .S0(clknet_1_0__leaf_net228),
    .S1(clknet_1_0__leaf_net968),
    .X(net236));
 sky130_fd_sc_hd__mux4_1 c242 (.A0(clknet_1_0__leaf_net227),
    .A1(net233),
    .A2(net224),
    .A3(clknet_1_0__leaf_net228),
    .S0(clknet_1_0__leaf_net926),
    .S1(net970),
    .X(net237));
 sky130_fd_sc_hd__mux4_1 c243 (.A0(net225),
    .A1(net233),
    .A2(clknet_1_1__leaf_net227),
    .A3(net884),
    .S0(clknet_1_0__leaf_net968),
    .S1(net973),
    .X(net238));
 sky130_fd_sc_hd__mux4_1 c244 (.A0(clknet_1_1__leaf_net226),
    .A1(net234),
    .A2(net224),
    .A3(clknet_1_1__leaf_net228),
    .S0(net971),
    .S1(net972),
    .X(net239));
 sky130_fd_sc_hd__mux4_1 c245 (.A0(net233),
    .A1(net225),
    .A2(clknet_1_0__leaf_net238),
    .A3(net971),
    .S0(net973),
    .S1(net975),
    .X(net240));
 sky130_fd_sc_hd__mux4_1 c246 (.A0(clknet_1_1__leaf_net238),
    .A1(clknet_1_1__leaf_net228),
    .A2(net234),
    .A3(net229),
    .S0(net972),
    .S1(net976),
    .X(net241));
 sky130_fd_sc_hd__mux4_1 c247 (.A0(net87),
    .A1(net233),
    .A2(net972),
    .A3(net975),
    .S0(net976),
    .S1(net977),
    .X(net242));
 sky130_fd_sc_hd__mux4_2 c248 (.A0(net225),
    .A1(net242),
    .A2(net224),
    .A3(net970),
    .S0(net974),
    .S1(net977),
    .X(net243));
 sky130_fd_sc_hd__mux4_1 c249 (.A0(net234),
    .A1(net243),
    .A2(clknet_1_1__leaf_net228),
    .A3(net974),
    .S0(net976),
    .S1(net977),
    .X(net244));
 sky130_fd_sc_hd__and3_1 c25 (.A(net1136),
    .B(net765),
    .C(net1138),
    .X(net0));
 sky130_fd_sc_hd__mux4_1 c250 (.A0(net243),
    .A1(clknet_1_1__leaf_net226),
    .A2(net809),
    .A3(net973),
    .S0(net976),
    .S1(net977),
    .X(net245));
 sky130_fd_sc_hd__mux4_1 c251 (.A0(net243),
    .A1(net866),
    .A2(net1149),
    .A3(net975),
    .S0(net976),
    .S1(net977),
    .X(net246));
 sky130_fd_sc_hd__and2_0 c252 (.A(clknet_1_1__leaf_net927),
    .B(net930),
    .X(net247));
 sky130_fd_sc_hd__and3_1 c253 (.A(clknet_1_1__leaf_net247),
    .B(clknet_1_1__leaf_net927),
    .C(net933),
    .X(net248));
 sky130_fd_sc_hd__and2_0 c254 (.A(clknet_1_0__leaf_net247),
    .B(clknet_1_1__leaf_net248),
    .X(net249));
 sky130_fd_sc_hd__sdfrtp_4 c255 (.CLK(clknet_leaf_10_clk),
    .D(clknet_1_0__leaf_net249),
    .RESET_B(clknet_1_0__leaf_net247),
    .SCD(clknet_1_0__leaf_net248),
    .SCE(clknet_1_1__leaf_net927),
    .Q(net250));
 sky130_fd_sc_hd__clkbuf_2 c256 (.A(net773),
    .X(net251));
 sky130_fd_sc_hd__or4bb_1 c257 (.A(net250),
    .B(clknet_1_0__leaf_net247),
    .C_N(net251),
    .D_N(clknet_1_0__leaf_net248),
    .X(net252));
 sky130_fd_sc_hd__buf_1 c258 (.A(net773),
    .X(net253));
 sky130_fd_sc_hd__sdfbbn_1 c259 (.CLK_N(clknet_leaf_11_clk),
    .D(net1260),
    .RESET_B(net253),
    .SCD(clknet_1_0__leaf_net248),
    .SCE(net250),
    .SET_B(clknet_1_1__leaf_net249),
    .Q(net255),
    .Q_N(net254));
 sky130_fd_sc_hd__or4bb_2 c26 (.A(net1139),
    .B(net631),
    .C_N(net1137),
    .D_N(net1136),
    .X(net1));
 sky130_fd_sc_hd__sdfbbn_1 c260 (.CLK_N(clknet_leaf_11_clk),
    .D(net1256),
    .RESET_B(clknet_1_1__leaf_net252),
    .SCD(net250),
    .SCE(clknet_1_0__leaf_net248),
    .SET_B(net1260),
    .Q(net257),
    .Q_N(net256));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(net251),
    .A1(clknet_1_0__leaf_net252),
    .A2(net256),
    .A3(clknet_1_1__leaf_net248),
    .S0(net250),
    .S1(net931),
    .X(net258));
 sky130_fd_sc_hd__mux4_1 c262 (.A0(clknet_1_0__leaf_net248),
    .A1(clknet_1_1__leaf_net249),
    .A2(net257),
    .A3(net253),
    .S0(net250),
    .S1(net251),
    .X(net259));
 sky130_fd_sc_hd__a2111o_1 c263 (.A1(net250),
    .A2(net251),
    .B1(net255),
    .C1(net256),
    .D1(clknet_1_1__leaf_net248),
    .X(net260));
 sky130_fd_sc_hd__mux4_1 c264 (.A0(net253),
    .A1(clknet_1_1__leaf_net260),
    .A2(net254),
    .A3(net250),
    .S0(net836),
    .S1(net979),
    .X(net261));
 sky130_fd_sc_hd__mux4_1 c265 (.A0(clknet_1_1__leaf_net247),
    .A1(net257),
    .A2(clknet_1_0__leaf_net260),
    .A3(clknet_1_1__leaf_net248),
    .S0(net253),
    .S1(net1202),
    .X(net262));
 sky130_fd_sc_hd__mux4_1 c266 (.A0(clknet_1_0__leaf_net260),
    .A1(net257),
    .A2(net250),
    .A3(net251),
    .S0(net1202),
    .S1(net981),
    .X(net263));
 sky130_fd_sc_hd__mux4_1 c267 (.A0(net257),
    .A1(net254),
    .A2(clknet_1_1__leaf_net260),
    .A3(net250),
    .S0(net1202),
    .S1(net984),
    .X(net264));
 sky130_fd_sc_hd__mux4_1 c268 (.A0(net1131),
    .A1(clknet_1_1__leaf_net260),
    .A2(net979),
    .A3(net1277),
    .S0(net984),
    .S1(net1244),
    .X(net265));
 sky130_fd_sc_hd__mux4_1 c269 (.A0(net253),
    .A1(net256),
    .A2(net836),
    .A3(net979),
    .S0(net981),
    .S1(net1244),
    .X(net266));
 sky130_fd_sc_hd__a2111o_4 c27 (.A1(net0),
    .A2(net811),
    .B1(net1135),
    .C1(net1),
    .D1(net1136),
    .X(net2));
 sky130_fd_sc_hd__mux4_1 c270 (.A0(net266),
    .A1(clknet_1_0__leaf_net260),
    .A2(net980),
    .A3(net981),
    .S0(net983),
    .S1(net985),
    .X(net267));
 sky130_fd_sc_hd__mux4_1 c271 (.A0(net266),
    .A1(clknet_1_0__leaf_net260),
    .A2(net868),
    .A3(net979),
    .S0(net984),
    .S1(net1244),
    .X(net268));
 sky130_fd_sc_hd__mux4_2 c272 (.A0(net117),
    .A1(net266),
    .A2(net856),
    .A3(net868),
    .S0(net983),
    .S1(net985),
    .X(net269));
 sky130_fd_sc_hd__and2_0 c273 (.A(net269),
    .B(net1202),
    .X(net270));
 sky130_fd_sc_hd__and2_1 c274 (.A(net154),
    .B(net269),
    .X(net271));
 sky130_fd_sc_hd__buf_1 c275 (.A(net763),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_2 c276 (.A(net867),
    .X(net273));
 sky130_fd_sc_hd__buf_1 c277 (.A(net763),
    .X(net274));
 sky130_fd_sc_hd__buf_1 c278 (.A(net793),
    .X(net275));
 sky130_fd_sc_hd__and3_1 c279 (.A(net272),
    .B(net273),
    .C(net1178),
    .X(net276));
 sky130_fd_sc_hd__and3_2 c28 (.A(net2),
    .B(net1136),
    .C(net1),
    .X(net3));
 sky130_fd_sc_hd__a2111o_1 c280 (.A1(net276),
    .A2(net1178),
    .B1(net272),
    .C1(net273),
    .D1(net1165),
    .X(net277));
 sky130_fd_sc_hd__buf_1 c281 (.A(clknet_1_0__leaf_net1128),
    .X(net278));
 sky130_fd_sc_hd__sdfbbp_1 c282 (.CLK(clknet_leaf_7_clk),
    .D(net271),
    .RESET_B(net1178),
    .SCD(net273),
    .SCE(net1257),
    .SET_B(net1225),
    .Q(net280),
    .Q_N(net279));
 sky130_fd_sc_hd__buf_1 c283 (.A(net1127),
    .X(net281));
 sky130_fd_sc_hd__mux4_1 c284 (.A0(net272),
    .A1(net1178),
    .A2(net1165),
    .A3(clknet_1_0__leaf_net278),
    .S0(net873),
    .S1(net1202),
    .X(net282));
 sky130_fd_sc_hd__sdfbbn_1 c285 (.CLK_N(clknet_leaf_7_clk),
    .D(net281),
    .RESET_B(net1178),
    .SCD(net1165),
    .SCE(net873),
    .SET_B(net1201),
    .Q(net284),
    .Q_N(net283));
 sky130_fd_sc_hd__mux4_1 c286 (.A0(net148),
    .A1(net275),
    .A2(net273),
    .A3(net274),
    .S0(net272),
    .S1(net1266),
    .X(net285));
 sky130_fd_sc_hd__mux4_1 c287 (.A0(net1165),
    .A1(net281),
    .A2(net272),
    .A3(net936),
    .S0(net1201),
    .S1(net1200),
    .X(net286));
 sky130_fd_sc_hd__mux4_1 c288 (.A0(net1165),
    .A1(net1178),
    .A2(net281),
    .A3(net1201),
    .S0(net1200),
    .S1(clknet_1_0__leaf_net988),
    .X(net287));
 sky130_fd_sc_hd__mux4_1 c289 (.A0(net1165),
    .A1(net153),
    .A2(net283),
    .A3(net1178),
    .S0(net1201),
    .S1(net1200),
    .X(net288));
 sky130_fd_sc_hd__sdfbbn_1 c29 (.CLK_N(clknet_leaf_2_clk),
    .D(net1138),
    .RESET_B(net3),
    .SCD(net1133),
    .SCE(net2),
    .SET_B(net1136),
    .Q(net5),
    .Q_N(net4));
 sky130_fd_sc_hd__mux4_1 c290 (.A0(net271),
    .A1(net1178),
    .A2(net273),
    .A3(net1201),
    .S0(net1200),
    .S1(clknet_1_1__leaf_net989),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 c291 (.A0(clknet_1_1__leaf_net278),
    .A1(net281),
    .A2(net269),
    .A3(net1200),
    .S0(clknet_1_1__leaf_net988),
    .S1(clknet_1_0__leaf_net990),
    .X(net290));
 sky130_fd_sc_hd__mux4_1 c292 (.A0(net284),
    .A1(clknet_1_1__leaf_net290),
    .A2(net1165),
    .A3(net1201),
    .S0(net1200),
    .S1(clknet_1_0__leaf_net989),
    .X(net291));
 sky130_fd_sc_hd__mux4_1 c293 (.A0(clknet_1_0__leaf_net290),
    .A1(net274),
    .A2(net273),
    .A3(net148),
    .S1(net992),
    .X(net292));
 sky130_fd_sc_hd__and2_0 c294 (.A(net1201),
    .B(net1200),
    .X(net293));
 sky130_fd_sc_hd__and2_1 c295 (.A(net1193),
    .B(net992),
    .X(net294));
 sky130_fd_sc_hd__and2_0 c296 (.A(net294),
    .B(net1193),
    .X(net295));
 sky130_fd_sc_hd__and2_1 c297 (.A(net1193),
    .B(net839),
    .X(net296));
 sky130_fd_sc_hd__and3_1 c298 (.A(net1193),
    .B(clknet_1_1__leaf_net948),
    .C(net1200),
    .X(net297));
 sky130_fd_sc_hd__or4bb_1 c299 (.A(net273),
    .B(clknet_1_0__leaf_net297),
    .C_N(net296),
    .D_N(net1193),
    .X(net298));
 sky130_fd_sc_hd__mux4_1 c30 (.A0(net754),
    .A1(net5),
    .A2(net0),
    .A3(net1137),
    .S0(net2),
    .S1(net3),
    .X(net6));
 sky130_fd_sc_hd__and3_1 c300 (.A(clknet_1_0__leaf_net297),
    .B(net1194),
    .C(net294),
    .X(net299));
 sky130_fd_sc_hd__a2111o_1 c301 (.A1(clknet_1_0__leaf_net298),
    .A2(net1193),
    .B1(net296),
    .C1(net295),
    .D1(net950),
    .X(net300));
 sky130_fd_sc_hd__mux4_1 c302 (.A0(clknet_1_0__leaf_net298),
    .A1(clknet_1_0__leaf_net297),
    .A2(net1194),
    .A3(net294),
    .S0(net296),
    .S1(net823),
    .X(net301));
 sky130_fd_sc_hd__sdfbbn_1 c303 (.CLK_N(clknet_leaf_6_clk),
    .D(clknet_1_1__leaf_net298),
    .RESET_B(net1194),
    .SCD(net296),
    .SCE(net294),
    .SET_B(net1246),
    .Q(net303),
    .Q_N(net302));
 sky130_fd_sc_hd__mux4_1 c304 (.A0(net303),
    .A1(clknet_1_1__leaf_net298),
    .A2(clknet_1_1__leaf_net297),
    .A3(net1193),
    .S0(clknet_1_1__leaf_net948),
    .S1(net993),
    .X(net304));
 sky130_fd_sc_hd__sdfbbp_1 c305 (.CLK(clknet_leaf_7_clk),
    .D(net299),
    .RESET_B(net294),
    .SCD(clknet_1_0__leaf_net298),
    .SCE(net1193),
    .SET_B(net993),
    .Q(net306),
    .Q_N(net305));
 sky130_fd_sc_hd__sdfbbn_1 c306 (.CLK_N(clknet_leaf_5_clk),
    .D(net295),
    .RESET_B(net1236),
    .SCD(net305),
    .SCE(net1193),
    .SET_B(net1229),
    .Q(net308),
    .Q_N(net307));
 sky130_fd_sc_hd__mux4_1 c307 (.A0(clknet_1_1__leaf_net297),
    .A1(net306),
    .A2(net302),
    .A3(net307),
    .S0(net294),
    .S1(net993),
    .X(net309));
 sky130_fd_sc_hd__sdfbbn_1 c308 (.CLK_N(clknet_leaf_5_clk),
    .D(net1262),
    .RESET_B(clknet_1_1__leaf_net298),
    .SCD(net305),
    .SCE(net1193),
    .SET_B(net1246),
    .Q(net311),
    .Q_N(net310));
 sky130_fd_sc_hd__mux4_2 c309 (.A0(net311),
    .A1(net302),
    .A2(net306),
    .A3(net1194),
    .S0(net823),
    .S1(net994),
    .X(net312));
 sky130_fd_sc_hd__mux4_1 c31 (.A0(net1),
    .A1(net9),
    .A2(net1137),
    .A3(net3),
    .S0(net4),
    .S1(net898),
    .X(net7));
 sky130_fd_sc_hd__mux4_1 c310 (.A0(net309),
    .A1(net312),
    .A2(net308),
    .A3(net305),
    .S0(net1194),
    .S1(net994),
    .X(net313));
 sky130_fd_sc_hd__mux4_2 c311 (.A0(net312),
    .A1(net310),
    .A2(net306),
    .A3(net307),
    .S0(net873),
    .S1(net994),
    .X(net314));
 sky130_fd_sc_hd__mux4_1 c312 (.A0(net311),
    .A1(net308),
    .A2(net303),
    .A3(net312),
    .S0(clknet_1_1__leaf_net297),
    .S1(net314),
    .X(net315));
 sky130_fd_sc_hd__mux4_1 c313 (.A0(net296),
    .A1(net306),
    .A2(net312),
    .A3(net310),
    .S0(net314),
    .S1(net307),
    .X(net316));
 sky130_fd_sc_hd__mux4_1 c314 (.A0(net296),
    .A1(net314),
    .A2(net311),
    .A3(net312),
    .S0(clknet_1_0__leaf_net891),
    .S1(net996),
    .X(net317));
 sky130_fd_sc_hd__or4bb_1 c315 (.A(clknet_1_0__leaf_net200),
    .B(net1195),
    .C_N(net182),
    .D_N(net996),
    .X(net318));
 sky130_fd_sc_hd__buf_1 c316 (.X(net319));
 sky130_fd_sc_hd__buf_2 c317 (.A(net764),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_2 c318 (.A(net1121),
    .X(net321));
 sky130_fd_sc_hd__sdfrtp_1 c319 (.CLK(clknet_leaf_42_clk),
    .D(net319),
    .RESET_B(clknet_1_1__leaf_net318),
    .SCD(net1195),
    .SCE(net320),
    .Q(net322));
 sky130_fd_sc_hd__mux4_1 c32 (.A0(net5),
    .A1(net2),
    .A2(net1),
    .A3(net3),
    .S0(net898),
    .S1(net899),
    .X(net8));
 sky130_fd_sc_hd__and3_1 c320 (.A(net321),
    .B(net306),
    .C(net320),
    .X(net323));
 sky130_fd_sc_hd__a2111o_1 c321 (.A1(net320),
    .A2(net1176),
    .B1(net321),
    .C1(clknet_1_0__leaf_net318),
    .D1(net322),
    .X(net324));
 sky130_fd_sc_hd__mux4_2 c322 (.A0(net182),
    .A1(net322),
    .A2(net321),
    .A3(net1176),
    .S0(net1200),
    .S1(net996),
    .X(net325));
 sky130_fd_sc_hd__buf_1 c323 (.A(net1122),
    .X(net326));
 sky130_fd_sc_hd__a2111o_2 c324 (.A1(net326),
    .A2(net321),
    .B1(net1177),
    .C1(net1195),
    .D1(net320),
    .X(net327));
 sky130_fd_sc_hd__sdfbbp_1 c325 (.CLK(clknet_leaf_43_clk),
    .D(clknet_1_0__leaf_net318),
    .RESET_B(net1250),
    .SCD(net320),
    .SCE(net327),
    .SET_B(net1176),
    .Q(net329),
    .Q_N(net328));
 sky130_fd_sc_hd__sdfbbn_1 c326 (.CLK_N(clknet_leaf_5_clk),
    .D(net329),
    .RESET_B(net1263),
    .SCD(net314),
    .SCE(net1176),
    .SET_B(net320),
    .Q(net331),
    .Q_N(net330));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(net327),
    .A1(net325),
    .A2(net326),
    .A3(net321),
    .S0(net1176),
    .S1(net881),
    .X(net332));
 sky130_fd_sc_hd__mux4_2 c328 (.A0(net331),
    .A1(net320),
    .A2(net328),
    .A3(net1176),
    .S0(net1195),
    .S1(net1201),
    .X(net333));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net333),
    .A1(net330),
    .A2(net327),
    .A3(net1176),
    .S0(net320),
    .S1(net328),
    .X(net334));
 sky130_fd_sc_hd__and2_0 c33 (.A(net1134),
    .B(net1133),
    .X(net9));
 sky130_fd_sc_hd__mux4_1 c330 (.A0(net332),
    .A1(net329),
    .A2(net333),
    .A3(net1177),
    .S0(net319),
    .S1(net334),
    .X(net335));
 sky130_fd_sc_hd__mux4_1 c331 (.A0(net334),
    .A1(net325),
    .A2(net322),
    .A3(net319),
    .S0(net333),
    .S1(net873),
    .X(net336));
 sky130_fd_sc_hd__mux4_1 c332 (.A0(net322),
    .A1(net333),
    .A2(net328),
    .A3(net1176),
    .S0(net881),
    .S1(net997),
    .X(net337));
 sky130_fd_sc_hd__mux4_1 c333 (.A0(net325),
    .A1(net329),
    .A2(clknet_1_0__leaf_net318),
    .A3(net321),
    .S0(net327),
    .S1(net997),
    .X(net338));
 sky130_fd_sc_hd__mux4_1 c334 (.A0(net333),
    .A1(net320),
    .A2(net319),
    .A3(net321),
    .S0(net995),
    .S1(net998),
    .X(net339));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(net337),
    .A1(net339),
    .A2(net329),
    .A3(net326),
    .S0(net997),
    .S1(net998),
    .X(net340));
 sky130_fd_sc_hd__or4bb_1 c336 (.A(net327),
    .B(net215),
    .C_N(clknet_1_1__leaf_net968),
    .D_N(clknet_1_1__leaf_net969),
    .X(net341));
 sky130_fd_sc_hd__sdfbbn_1 c337 (.CLK_N(clknet_leaf_41_clk),
    .D(clknet_1_0__leaf_net341),
    .RESET_B(net1177),
    .SCD(net214),
    .SCE(clknet_1_1__leaf_net968),
    .SET_B(clknet_1_1__leaf_net969),
    .Q(net343),
    .Q_N(net342));
 sky130_fd_sc_hd__sdfsbp_1 c338 (.CLK(clknet_leaf_41_clk),
    .D(net343),
    .SCD(net1177),
    .SCE(clknet_1_0__leaf_net341),
    .SET_B(clknet_1_1__leaf_net968),
    .Q(net345),
    .Q_N(net344));
 sky130_fd_sc_hd__sdfbbp_1 c339 (.CLK(clknet_leaf_41_clk),
    .D(net1273),
    .RESET_B(net1177),
    .SCD(net215),
    .SCE(net342),
    .SET_B(clknet_1_0__leaf_net341),
    .Q(net347),
    .Q_N(net346));
 sky130_fd_sc_hd__mux4_1 c34 (.A0(net3),
    .A1(net1144),
    .A2(net1129),
    .A3(net5),
    .S0(net2),
    .S1(net897),
    .X(net10));
 sky130_fd_sc_hd__sdfbbn_1 c340 (.CLK_N(clknet_leaf_41_clk),
    .D(net347),
    .RESET_B(net1248),
    .SCD(net325),
    .SCE(clknet_1_0__leaf_net341),
    .SET_B(net1177),
    .Q(net349),
    .Q_N(net348));
 sky130_fd_sc_hd__sdfbbn_1 c341 (.CLK_N(clknet_leaf_41_clk),
    .D(net1268),
    .RESET_B(clknet_1_1__leaf_net341),
    .SCD(net1248),
    .SCE(net346),
    .SET_B(net1177),
    .Q(net351),
    .Q_N(net350));
 sky130_fd_sc_hd__sdfbbp_1 c342 (.CLK(clknet_leaf_40_clk),
    .D(net349),
    .RESET_B(clknet_1_0__leaf_net341),
    .SCD(net351),
    .SCE(net342),
    .SET_B(net344),
    .Q(net353),
    .Q_N(net352));
 sky130_fd_sc_hd__mux4_1 c343 (.A0(net353),
    .A1(net349),
    .A2(net351),
    .A3(net346),
    .S0(clknet_1_1__leaf_net341),
    .S1(net342),
    .X(net354));
 sky130_fd_sc_hd__sdfbbn_1 c344 (.CLK_N(clknet_leaf_40_clk),
    .D(net1264),
    .RESET_B(net352),
    .SCD(net1171),
    .SCE(clknet_1_0__leaf_net341),
    .SET_B(net1199),
    .Q(net356),
    .Q_N(net355));
 sky130_fd_sc_hd__mux4_1 c345 (.A0(net343),
    .A1(net350),
    .A2(net355),
    .A3(clknet_1_1__leaf_net341),
    .S0(net999),
    .S1(net1199),
    .X(net357));
 sky130_fd_sc_hd__mux4_1 c346 (.A0(net353),
    .A1(net356),
    .A2(net348),
    .A3(net350),
    .S0(net1199),
    .S1(net1001),
    .X(net358));
 sky130_fd_sc_hd__mux4_2 c347 (.A0(net358),
    .A1(net344),
    .A2(net356),
    .A3(net350),
    .S0(net1199),
    .S1(net1001),
    .X(net359));
 sky130_fd_sc_hd__mux4_1 c348 (.A0(net358),
    .A1(net359),
    .A2(net356),
    .A3(net348),
    .S0(net342),
    .S1(net350),
    .X(net360));
 sky130_fd_sc_hd__mux4_1 c349 (.A0(net360),
    .A1(net351),
    .A2(net359),
    .A3(net348),
    .S0(net1199),
    .S1(net1001),
    .X(net361));
 sky130_fd_sc_hd__mux4_1 c35 (.A0(net1142),
    .A1(net4),
    .A2(net2),
    .A3(net898),
    .S0(net900),
    .S1(net901),
    .X(net11));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(net349),
    .A1(net355),
    .A2(net359),
    .A3(clknet_1_1__leaf_net341),
    .S0(net1199),
    .S1(net1003),
    .X(net362));
 sky130_fd_sc_hd__mux4_2 c351 (.A0(net356),
    .A1(net359),
    .A2(net358),
    .A3(net1199),
    .S0(net1003),
    .S1(net1004),
    .X(net363));
 sky130_fd_sc_hd__mux4_1 c352 (.A0(net363),
    .A1(net360),
    .A2(net359),
    .A3(net355),
    .S0(net1003),
    .S1(net1271),
    .X(net364));
 sky130_fd_sc_hd__mux4_1 c353 (.A0(net363),
    .A1(net327),
    .A2(net359),
    .A3(net1002),
    .S0(net1285),
    .S1(net1280),
    .X(net365));
 sky130_fd_sc_hd__mux4_1 c354 (.A0(net345),
    .A1(net358),
    .A2(net363),
    .A3(net1004),
    .S0(net1006),
    .S1(net1223),
    .X(net366));
 sky130_fd_sc_hd__mux4_1 c355 (.A0(clknet_1_1__leaf_net341),
    .A1(net360),
    .A2(net363),
    .S0(net1001),
    .S1(net1007),
    .X(net367));
 sky130_fd_sc_hd__sdfbbn_1 c356 (.CLK_N(clknet_leaf_38_clk),
    .D(net363),
    .RESET_B(net812),
    .SCD(net1002),
    .SCE(net1006),
    .SET_B(net1007),
    .Q(net369),
    .Q_N(net368));
 sky130_fd_sc_hd__and3_1 c357 (.A(net369),
    .B(net325),
    .C(net810),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_2 c358 (.A(net1123),
    .X(net371));
 sky130_fd_sc_hd__and2_1 c359 (.A(net369),
    .B(net371),
    .X(net372));
 sky130_fd_sc_hd__mux4_1 c36 (.A0(net9),
    .A1(net781),
    .A2(net2),
    .A3(net4),
    .S0(net898),
    .S1(net901),
    .X(net12));
 sky130_fd_sc_hd__a2111o_2 c360 (.A1(net1175),
    .A2(net346),
    .B1(net369),
    .C1(net1230),
    .D1(net1218),
    .X(net373));
 sky130_fd_sc_hd__a2111o_1 c361 (.A1(net371),
    .A2(net1175),
    .B1(net373),
    .C1(net368),
    .D1(net1000),
    .X(net374));
 sky130_fd_sc_hd__a2111o_1 c362 (.A1(net243),
    .A2(net1175),
    .B1(net373),
    .C1(net1164),
    .D1(net1230),
    .X(net375));
 sky130_fd_sc_hd__mux4_1 c363 (.A0(net224),
    .A1(net1164),
    .A2(net371),
    .A3(net368),
    .S0(net1175),
    .S1(net373),
    .X(net376));
 sky130_fd_sc_hd__mux4_1 c364 (.A0(net373),
    .A1(net1175),
    .A2(net1164),
    .A3(net368),
    .S0(net371),
    .S1(net1008),
    .X(net377));
 sky130_fd_sc_hd__mux4_1 c365 (.A0(clknet_1_1__leaf_net105),
    .A1(net373),
    .A2(net1164),
    .A3(net1175),
    .S0(net1008),
    .S1(clknet_1_0__leaf_net1009),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 c366 (.A0(net371),
    .A1(net1175),
    .A2(net1164),
    .A3(net815),
    .S0(net1008),
    .S1(clknet_1_0__leaf_net1009),
    .X(net379));
 sky130_fd_sc_hd__mux4_1 c367 (.A0(net1175),
    .A1(net1164),
    .A2(net815),
    .A3(net1008),
    .S0(clknet_1_0__leaf_net1009),
    .S1(clknet_1_0__leaf_net1011),
    .X(net380));
 sky130_fd_sc_hd__mux4_1 c368 (.A0(net369),
    .A1(net1175),
    .A2(net1008),
    .A3(clknet_1_0__leaf_net1009),
    .S0(clknet_1_0__leaf_net1010),
    .S1(net1013),
    .X(net381));
 sky130_fd_sc_hd__mux4_1 c369 (.A0(net1164),
    .A1(clknet_1_0__leaf_net381),
    .A2(net1175),
    .A3(net1008),
    .S0(clknet_1_1__leaf_net1009),
    .S1(net1013),
    .X(net382));
 sky130_fd_sc_hd__mux4_1 c37 (.A0(net12),
    .A1(net11),
    .A2(net3),
    .A3(net897),
    .S0(net900),
    .S1(net901),
    .X(net13));
 sky130_fd_sc_hd__mux4_1 c370 (.A0(net1164),
    .A1(net372),
    .A2(net1008),
    .A3(clknet_1_1__leaf_net1009),
    .S0(net1013),
    .S1(net1015),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(net370),
    .A1(net373),
    .A2(clknet_1_0__leaf_net1009),
    .A3(clknet_1_1__leaf_net1011),
    .S0(net1012),
    .S1(net1014),
    .X(net384));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(clknet_1_0__leaf_net381),
    .A1(net1008),
    .A2(net1012),
    .A3(net1015),
    .S0(net1016),
    .S1(net1018),
    .X(net385));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net374),
    .A1(clknet_1_0__leaf_net385),
    .A2(net1008),
    .A3(clknet_1_1__leaf_net1009),
    .S0(clknet_1_1__leaf_net1010),
    .S1(net1015),
    .X(net386));
 sky130_fd_sc_hd__mux4_1 c374 (.A0(clknet_1_1__leaf_net381),
    .A1(clknet_1_1__leaf_net385),
    .A2(net1164),
    .A3(net372),
    .S0(clknet_1_1__leaf_net1009),
    .S1(net1019),
    .X(net387));
 sky130_fd_sc_hd__mux4_1 c375 (.A0(clknet_1_1__leaf_net385),
    .A1(clknet_1_1__leaf_net381),
    .A2(net893),
    .A3(clknet_1_1__leaf_net1009),
    .S0(net1014),
    .S1(net1017),
    .X(net388));
 sky130_fd_sc_hd__mux4_1 c376 (.A0(clknet_1_1__leaf_net381),
    .A1(clknet_1_1__leaf_net385),
    .A2(net861),
    .A3(net1008),
    .S0(net1018),
    .S1(net1019),
    .X(net389));
 sky130_fd_sc_hd__mux4_1 c377 (.A0(net371),
    .A1(clknet_1_0__leaf_net385),
    .A2(net1164),
    .A3(net815),
    .S0(net861),
    .S1(net893),
    .X(net390));
 sky130_fd_sc_hd__and2_0 c378 (.A(net1202),
    .B(net982),
    .X(net391));
 sky130_fd_sc_hd__and2_0 c379 (.A(net391),
    .B(net1202),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c38 (.A0(net1137),
    .A1(net2),
    .A2(net5),
    .A3(net897),
    .S0(net901),
    .S1(net902),
    .X(net14));
 sky130_fd_sc_hd__and2_0 c380 (.A(net392),
    .B(net269),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_1 c381 (.X(net394));
 sky130_fd_sc_hd__and2_1 c382 (.A(net269),
    .B(net1225),
    .X(net395));
 sky130_fd_sc_hd__buf_1 c383 (.A(net779),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_1 c384 (.A(net786),
    .X(net397));
 sky130_fd_sc_hd__sdfsbp_1 c385 (.CLK(clknet_leaf_12_clk),
    .D(net1237),
    .SCD(net1210),
    .SCE(net1191),
    .SET_B(net395),
    .Q(net399),
    .Q_N(net398));
 sky130_fd_sc_hd__or4bb_4 c386 (.A(net1210),
    .B(net1191),
    .C_N(net1202),
    .D_N(net982),
    .X(net400));
 sky130_fd_sc_hd__sdfbbp_1 c387 (.CLK(clknet_leaf_12_clk),
    .D(net400),
    .RESET_B(net1191),
    .SCD(net395),
    .SCE(net1210),
    .SET_B(net1220),
    .Q(net402),
    .Q_N(net401));
 sky130_fd_sc_hd__a2111o_1 c388 (.A1(net1210),
    .A2(net399),
    .B1(net402),
    .C1(net400),
    .D1(net1191),
    .X(net403));
 sky130_fd_sc_hd__mux4_2 c389 (.A0(net392),
    .A1(net403),
    .A2(net1210),
    .A3(net402),
    .S0(net1191),
    .S1(net1202),
    .X(net404));
 sky130_fd_sc_hd__mux4_1 c39 (.A0(net3),
    .A1(net1136),
    .A2(net2),
    .A3(clknet_1_0__leaf_net855),
    .S0(net901),
    .S1(net902),
    .X(net15));
 sky130_fd_sc_hd__mux4_1 c390 (.A0(net403),
    .A1(net400),
    .A2(net404),
    .A3(net401),
    .S0(net1191),
    .S1(net1210),
    .X(net405));
 sky130_fd_sc_hd__mux4_1 c391 (.A0(net395),
    .A1(net403),
    .A2(net402),
    .A3(net1191),
    .S0(net400),
    .S1(net1210),
    .X(net406));
 sky130_fd_sc_hd__mux4_1 c392 (.A0(net402),
    .A1(net400),
    .A2(net403),
    .A3(net1191),
    .S0(net1210),
    .S1(net840),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net402),
    .A1(net400),
    .A2(net403),
    .A3(net1191),
    .S0(net1210),
    .S1(net840),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c394 (.A0(net407),
    .A1(net400),
    .A2(net403),
    .A3(net396),
    .S0(net401),
    .S1(net404),
    .X(net409));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net404),
    .A1(net407),
    .A2(net396),
    .A3(net401),
    .S0(net400),
    .S1(net1021),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 c396 (.A0(net408),
    .A1(net400),
    .A2(net1192),
    .A3(net401),
    .S0(net1021),
    .S1(net1261),
    .X(net411));
 sky130_fd_sc_hd__mux4_1 c397 (.A0(net408),
    .A1(net404),
    .A2(net840),
    .A3(net1021),
    .S0(net1261),
    .S1(net1023),
    .X(net412));
 sky130_fd_sc_hd__mux4_1 c398 (.A0(net391),
    .A1(net400),
    .A2(net840),
    .A3(net1021),
    .S0(net1024),
    .S1(net1026),
    .X(net413));
 sky130_fd_sc_hd__and2_0 c399 (.A(net937),
    .B(net1239),
    .X(net414));
 sky130_fd_sc_hd__mux4_1 c40 (.A0(net14),
    .A1(net1146),
    .A2(net811),
    .A3(net5),
    .S0(clknet_1_0__leaf_net855),
    .S1(net902),
    .X(net16));
 sky130_fd_sc_hd__and2_1 c400 (.A(net1201),
    .B(net992),
    .X(net415));
 sky130_fd_sc_hd__and2_2 c401 (.A(net987),
    .B(net991),
    .X(net416));
 sky130_fd_sc_hd__and3_1 c402 (.A(net416),
    .B(net415),
    .C(clknet_1_1__leaf_net990),
    .X(net417));
 sky130_fd_sc_hd__and3_1 c403 (.A(clknet_1_0__leaf_net417),
    .B(net415),
    .C(net416),
    .X(net418));
 sky130_fd_sc_hd__sdfbbn_1 c404 (.CLK_N(clknet_leaf_15_clk),
    .D(clknet_1_0__leaf_net418),
    .RESET_B(net414),
    .SCD(net416),
    .SCE(net279),
    .SET_B(net415),
    .Q(net420),
    .Q_N(net419));
 sky130_fd_sc_hd__buf_1 c405 (.A(net790),
    .X(net421));
 sky130_fd_sc_hd__sdfbbn_1 c406 (.CLK_N(clknet_leaf_15_clk),
    .D(net414),
    .RESET_B(net415),
    .SCD(clknet_1_0__leaf_net418),
    .SCE(net420),
    .SET_B(net1190),
    .Q(net423),
    .Q_N(net422));
 sky130_fd_sc_hd__a2111o_1 c407 (.A1(net415),
    .A2(net423),
    .B1(net420),
    .C1(net1190),
    .D1(net416),
    .X(net424));
 sky130_fd_sc_hd__a2111o_1 c408 (.A1(net1190),
    .A2(net420),
    .B1(net422),
    .C1(net416),
    .D1(net1247),
    .X(net425));
 sky130_fd_sc_hd__a2111o_2 c409 (.A1(net423),
    .A2(net1190),
    .B1(net425),
    .C1(net416),
    .D1(net419),
    .X(net426));
 sky130_fd_sc_hd__mux4_1 c41 (.A0(net2),
    .A1(net12),
    .A2(net4),
    .A3(net3),
    .S0(net880),
    .S1(net902),
    .X(net17));
 sky130_fd_sc_hd__sdfbbp_1 c410 (.CLK(clknet_leaf_15_clk),
    .D(clknet_1_0__leaf_net417),
    .RESET_B(net420),
    .SCD(net1190),
    .SCE(net426),
    .SET_B(net425),
    .Q(net428),
    .Q_N(net427));
 sky130_fd_sc_hd__mux4_1 c411 (.A0(net420),
    .A1(net416),
    .A2(net425),
    .A3(net426),
    .S0(net427),
    .S1(net421),
    .X(net429));
 sky130_fd_sc_hd__sdfbbn_1 c412 (.CLK_N(clknet_leaf_7_clk),
    .D(net428),
    .RESET_B(net426),
    .SCD(net1190),
    .SCE(net419),
    .SET_B(net1201),
    .Q(net431),
    .Q_N(net430));
 sky130_fd_sc_hd__mux4_1 c413 (.A0(net425),
    .A1(net426),
    .A2(net427),
    .A3(net419),
    .S0(net1190),
    .S1(net422),
    .X(net432));
 sky130_fd_sc_hd__mux4_1 c414 (.A0(net416),
    .A1(net428),
    .A2(net423),
    .A3(net426),
    .S0(net1190),
    .S1(net1265),
    .X(net433));
 sky130_fd_sc_hd__mux4_1 c415 (.A0(net431),
    .A1(net415),
    .A2(net1190),
    .A3(net426),
    .S0(net1282),
    .S1(net422),
    .X(net434));
 sky130_fd_sc_hd__sdfbbn_1 c416 (.CLK_N(clknet_leaf_16_clk),
    .D(net428),
    .RESET_B(net426),
    .SCD(net1190),
    .SCE(net1027),
    .SET_B(net1028),
    .Q(net436),
    .Q_N(net435));
 sky130_fd_sc_hd__mux4_1 c417 (.A0(net426),
    .A1(clknet_1_1__leaf_net417),
    .A2(net419),
    .A3(net422),
    .S0(net421),
    .S1(net825),
    .X(net437));
 sky130_fd_sc_hd__mux4_1 c418 (.A0(net424),
    .A1(net430),
    .A2(net423),
    .A3(net427),
    .S0(net426),
    .X(net438));
 sky130_fd_sc_hd__mux4_1 c419 (.A0(net428),
    .A1(net423),
    .A2(net435),
    .A3(net426),
    .S0(net871),
    .S1(net1028),
    .X(net439));
 sky130_fd_sc_hd__and3_1 c42 (.A(net794),
    .B(net811),
    .C(net1204),
    .X(net18));
 sky130_fd_sc_hd__buf_1 c420 (.A(net831),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_1 c421 (.A(net830),
    .X(net441));
 sky130_fd_sc_hd__and2_1 c422 (.A(net1186),
    .B(net1188),
    .X(net442));
 sky130_fd_sc_hd__and3_1 c423 (.A(net1186),
    .B(net1188),
    .C(net996),
    .X(net443));
 sky130_fd_sc_hd__and3_1 c424 (.A(net1188),
    .B(net1186),
    .C(net995),
    .X(net444));
 sky130_fd_sc_hd__and3_1 c425 (.A(net1188),
    .B(net444),
    .C(net1186),
    .X(net445));
 sky130_fd_sc_hd__and3_1 c426 (.A(net1189),
    .B(net442),
    .C(net857),
    .X(net446));
 sky130_fd_sc_hd__or4bb_1 c427 (.A(net445),
    .B(net1186),
    .C_N(net446),
    .D_N(net1189),
    .X(net447));
 sky130_fd_sc_hd__mux4_2 c428 (.A0(net442),
    .A1(net444),
    .A2(net446),
    .A3(net1187),
    .S0(net1188),
    .S1(net445),
    .X(net448));
 sky130_fd_sc_hd__sdfbbp_1 c429 (.CLK(clknet_leaf_16_clk),
    .D(net446),
    .RESET_B(net444),
    .SCD(net448),
    .SCE(net1187),
    .SET_B(net1188),
    .Q(net450),
    .Q_N(net449));
 sky130_fd_sc_hd__and2_1 c43 (.A(net18),
    .B(net1203),
    .X(net19));
 sky130_fd_sc_hd__mux4_1 c430 (.A0(net450),
    .A1(net1189),
    .A2(net305),
    .A3(net1187),
    .S0(net448),
    .S1(net1281),
    .X(net451));
 sky130_fd_sc_hd__mux4_1 c431 (.A0(net306),
    .A1(net445),
    .A2(net1186),
    .A3(net1188),
    .S0(net448),
    .S1(net1198),
    .X(net452));
 sky130_fd_sc_hd__mux4_1 c432 (.A0(net448),
    .A1(net1187),
    .A2(net305),
    .A3(net1189),
    .S0(net1198),
    .S1(clknet_1_1__leaf_net1030),
    .X(net453));
 sky130_fd_sc_hd__mux4_1 c433 (.A0(net314),
    .A1(net445),
    .A2(net1186),
    .A3(net1188),
    .S0(net1198),
    .S1(clknet_1_0__leaf_net1031),
    .X(net454));
 sky130_fd_sc_hd__mux4_1 c434 (.A0(net450),
    .A1(net1187),
    .A2(net1189),
    .A3(clknet_1_0__leaf_net1030),
    .S0(clknet_1_0__leaf_net1031),
    .S1(clknet_1_1__leaf_net1032),
    .X(net455));
 sky130_fd_sc_hd__mux4_1 c435 (.A0(net447),
    .A1(net1188),
    .A2(net1186),
    .A3(net1198),
    .S0(clknet_1_0__leaf_net1031),
    .S1(clknet_1_0__leaf_net1032),
    .X(net456));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net449),
    .A1(net1187),
    .A2(net1198),
    .A3(clknet_1_0__leaf_net1030),
    .S0(clknet_1_1__leaf_net1031),
    .S1(net1034),
    .X(net457));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(net455),
    .A1(clknet_1_1__leaf_net457),
    .A2(net1186),
    .A3(net1198),
    .S0(clknet_1_1__leaf_net1031),
    .S1(net1034),
    .X(net458));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(clknet_1_0__leaf_net458),
    .A1(clknet_1_0__leaf_net457),
    .A2(net1186),
    .A3(net442),
    .S0(clknet_1_1__leaf_net1031),
    .S1(clknet_1_0__leaf_net1032),
    .X(net459));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net443),
    .A1(clknet_1_0__leaf_net457),
    .A2(net448),
    .A3(clknet_1_0__leaf_net458),
    .S0(clknet_1_0__leaf_net1031),
    .S1(net1033),
    .X(net460));
 sky130_fd_sc_hd__and2_1 c44 (.A(net18),
    .B(net1204),
    .X(net20));
 sky130_fd_sc_hd__mux4_1 c440 (.A0(net459),
    .A1(clknet_1_1__leaf_net458),
    .A2(clknet_1_1__leaf_net457),
    .A3(net831),
    .S0(net1198),
    .S1(clknet_1_1__leaf_net1031),
    .X(net461));
 sky130_fd_sc_hd__and2_1 c441 (.A(net999),
    .B(net1036),
    .X(net462));
 sky130_fd_sc_hd__and2_1 c442 (.A(net462),
    .B(net1198),
    .X(net463));
 sky130_fd_sc_hd__and3_1 c443 (.A(net463),
    .B(net325),
    .C(net1176),
    .X(net464));
 sky130_fd_sc_hd__buf_1 c444 (.A(clknet_1_1__leaf_net890),
    .X(net465));
 sky130_fd_sc_hd__sdfstp_1 c445 (.CLK(clknet_leaf_42_clk),
    .D(net463),
    .SCD(clknet_1_0__leaf_net465),
    .SCE(net1163),
    .SET_B(net1036),
    .Q(net466));
 sky130_fd_sc_hd__sdfbbn_1 c446 (.CLK_N(clknet_leaf_42_clk),
    .D(clknet_1_1__leaf_net181),
    .RESET_B(net466),
    .SCD(clknet_1_0__leaf_net465),
    .SCE(net1163),
    .SET_B(net1242),
    .Q(net468),
    .Q_N(net467));
 sky130_fd_sc_hd__buf_1 c447 (.A(clknet_1_1__leaf_net890),
    .X(net469));
 sky130_fd_sc_hd__mux4_1 c448 (.A0(clknet_1_0__leaf_net465),
    .A1(net466),
    .A2(net1163),
    .A3(net462),
    .S0(net999),
    .S1(net1198),
    .X(net470));
 sky130_fd_sc_hd__sdfbbn_1 c449 (.CLK_N(clknet_leaf_42_clk),
    .D(net466),
    .RESET_B(net1254),
    .SCD(net1163),
    .SCE(clknet_1_0__leaf_net465),
    .SET_B(net1242),
    .Q(net472),
    .Q_N(net471));
 sky130_fd_sc_hd__and3_1 c45 (.A(net1174),
    .B(net19),
    .C(net1203),
    .X(net21));
 sky130_fd_sc_hd__sdfbbp_1 c450 (.CLK(clknet_leaf_42_clk),
    .D(net1163),
    .RESET_B(clknet_1_1__leaf_net465),
    .SCD(net471),
    .SCE(net1279),
    .SET_B(net1038),
    .Q(net474),
    .Q_N(net473));
 sky130_fd_sc_hd__mux4_1 c451 (.A0(net474),
    .A1(net466),
    .A2(clknet_1_1__leaf_net465),
    .A3(net471),
    .S0(net1163),
    .S1(net1177),
    .X(net475));
 sky130_fd_sc_hd__sdfbbn_1 c452 (.CLK_N(clknet_leaf_29_clk),
    .D(net1258),
    .RESET_B(net474),
    .SCD(net1163),
    .SCE(clknet_1_0__leaf_net465),
    .SET_B(net1251),
    .Q(net477),
    .Q_N(net476));
 sky130_fd_sc_hd__mux4_1 c453 (.A0(net477),
    .A1(clknet_1_0__leaf_net469),
    .A2(net472),
    .A3(net473),
    .S0(clknet_1_1__leaf_net465),
    .S1(net1163),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c454 (.A0(clknet_1_0__leaf_net469),
    .A1(net477),
    .A2(net474),
    .A3(net472),
    .S0(net1036),
    .S1(net1040),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c455 (.A0(net280),
    .A1(clknet_1_1__leaf_net479),
    .A2(net464),
    .A3(net473),
    .S0(net1039),
    .S1(net1040),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(clknet_1_1__leaf_net465),
    .A1(net474),
    .A2(net476),
    .A3(net1163),
    .S0(net1040),
    .S1(net1041),
    .X(net481));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(clknet_1_0__leaf_net479),
    .A1(net467),
    .A2(net473),
    .A3(net879),
    .S0(net1039),
    .S1(net1040),
    .X(net482));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(clknet_1_1__leaf_net482),
    .A1(clknet_1_1__leaf_net469),
    .A2(clknet_1_0__leaf_net479),
    .A3(net473),
    .S0(net1040),
    .S1(net1041),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net468),
    .A1(clknet_1_0__leaf_net483),
    .A2(clknet_1_0__leaf_net482),
    .A3(net471),
    .S0(net1039),
    .S1(net1041),
    .X(net484));
 sky130_fd_sc_hd__clkbuf_1 c46 (.A(net865),
    .X(net22));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net462),
    .A1(net468),
    .A2(clknet_1_0__leaf_net483),
    .A3(net1149),
    .S0(net999),
    .S1(net1037),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(clknet_1_1__leaf_net483),
    .A1(clknet_1_0__leaf_net482),
    .A2(net1149),
    .A3(net1040),
    .S0(net1041),
    .S1(net1197),
    .X(net486));
 sky130_fd_sc_hd__and3_1 c462 (.A(net347),
    .B(clknet_1_1__leaf_net968),
    .C(net1199),
    .X(net487));
 sky130_fd_sc_hd__and3_1 c463 (.A(clknet_1_0__leaf_net487),
    .B(net346),
    .C(net1197),
    .X(net488));
 sky130_fd_sc_hd__and3_1 c464 (.A(clknet_1_0__leaf_net488),
    .B(clknet_1_0__leaf_net487),
    .C(net323),
    .X(net489));
 sky130_fd_sc_hd__sdfbbn_1 c465 (.CLK_N(clknet_leaf_30_clk),
    .D(net359),
    .RESET_B(clknet_1_1__leaf_net489),
    .SCD(clknet_1_0__leaf_net488),
    .SCE(net1035),
    .SET_B(net1197),
    .Q(net491),
    .Q_N(net490));
 sky130_fd_sc_hd__a2111o_1 c466 (.A1(net491),
    .A2(clknet_1_1__leaf_net487),
    .B1(clknet_1_0__leaf_net488),
    .C1(net879),
    .D1(net1199),
    .X(net492));
 sky130_fd_sc_hd__mux4_1 c467 (.A0(clknet_1_0__leaf_net489),
    .A1(clknet_1_1__leaf_net200),
    .A2(net490),
    .A3(net359),
    .S0(clknet_1_0__leaf_net488),
    .S1(clknet_1_0__leaf_net487),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c468 (.A0(clknet_1_0__leaf_net488),
    .A1(clknet_1_1__leaf_net492),
    .A2(net490),
    .A3(clknet_1_1__leaf_net487),
    .S0(net1035),
    .S1(net1043),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c469 (.A0(net491),
    .A1(clknet_1_1__leaf_net492),
    .A2(clknet_1_1__leaf_net489),
    .A3(clknet_1_1__leaf_net487),
    .S0(clknet_1_0__leaf_net488),
    .S1(net1043),
    .X(net495));
 sky130_fd_sc_hd__clkbuf_1 c47 (.A(net865),
    .X(net23));
 sky130_fd_sc_hd__mux4_1 c470 (.A0(clknet_1_1__leaf_net488),
    .A1(clknet_1_0__leaf_net492),
    .A2(clknet_1_0__leaf_net487),
    .A3(net1199),
    .S0(net1043),
    .S1(net1044),
    .X(net496));
 sky130_fd_sc_hd__a2111o_1 c471 (.A1(clknet_1_1__leaf_net487),
    .A2(clknet_1_1__leaf_net488),
    .B1(clknet_1_1__leaf_net492),
    .D1(net1046),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c472 (.A0(clknet_1_0__leaf_net489),
    .A1(clknet_1_1__leaf_net488),
    .A2(clknet_1_0__leaf_net487),
    .A3(clknet_1_0__leaf_net492),
    .S0(net1043),
    .S1(net1046),
    .X(net498));
 sky130_fd_sc_hd__a2111o_1 c473 (.A1(clknet_1_1__leaf_net488),
    .A2(clknet_1_0__leaf_net487),
    .B1(net835),
    .C1(net1000),
    .D1(net1047),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c474 (.A0(clknet_1_1__leaf_net488),
    .A1(clknet_1_0__leaf_net489),
    .A2(clknet_1_0__leaf_net487),
    .A3(net1044),
    .S0(net1046),
    .S1(net1048),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c475 (.A0(clknet_1_1__leaf_net489),
    .A1(clknet_1_1__leaf_net487),
    .A2(net490),
    .A3(net834),
    .S0(net1045),
    .S1(net1047),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(clknet_1_0__leaf_net492),
    .A1(clknet_1_0__leaf_net499),
    .A2(clknet_1_1__leaf_net488),
    .A3(clknet_1_0__leaf_net487),
    .S0(net1046),
    .S1(net1156),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c477 (.A0(net347),
    .A1(clknet_1_1__leaf_net488),
    .A2(clknet_1_0__leaf_net487),
    .A3(net1047),
    .S0(net1048),
    .S1(net1156),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(clknet_1_1__leaf_net499),
    .A1(clknet_1_0__leaf_net503),
    .A2(net1043),
    .A3(net1048),
    .S0(net1049),
    .S1(net1156),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(clknet_1_0__leaf_net503),
    .A1(clknet_1_1__leaf_net487),
    .A2(net1197),
    .A3(net1045),
    .S0(net1048),
    .S1(net1156),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_1 c48 (.A(net1127),
    .X(net24));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(clknet_1_1__leaf_net503),
    .A1(net1043),
    .A2(net1044),
    .A3(net1049),
    .S0(clknet_1_1__leaf_net1051),
    .S1(clknet_1_1__leaf_net1052),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(clknet_1_1__leaf_net487),
    .A1(net491),
    .A2(clknet_1_0__leaf_net892),
    .A3(net1045),
    .S0(net1048),
    .S1(clknet_1_0__leaf_net1051),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(clknet_1_1__leaf_net503),
    .A1(clknet_1_0__leaf_net892),
    .A2(net1197),
    .A3(net1047),
    .S0(net1048),
    .S1(clknet_1_0__leaf_net1052),
    .X(net508));
 sky130_fd_sc_hd__and2_0 c483 (.A(clknet_1_0__leaf_net507),
    .B(net1020),
    .X(net1150));
 sky130_fd_sc_hd__buf_1 c484 (.A(net772),
    .X(net509));
 sky130_fd_sc_hd__buf_1 c485 (.A(net772),
    .X(net510));
 sky130_fd_sc_hd__and3_1 c486 (.A(net509),
    .B(clknet_1_0__leaf_net507),
    .C(net510),
    .X(net1160));
 sky130_fd_sc_hd__buf_1 c487 (.A(net1124),
    .X(net1161));
 sky130_fd_sc_hd__sdfbbp_1 c488 (.CLK(clknet_leaf_34_clk),
    .D(net510),
    .RESET_B(net1161),
    .SCD(clknet_1_0__leaf_net1160),
    .SCE(clknet_1_0__leaf_net1150),
    .SET_B(clknet_1_0__leaf_net1050),
    .Q(net512),
    .Q_N(net511));
 sky130_fd_sc_hd__buf_1 c489 (.A(net894),
    .X(net1162));
 sky130_fd_sc_hd__buf_2 c49 (.A(net1126),
    .X(net25));
 sky130_fd_sc_hd__sdfbbn_1 c490 (.CLK_N(clknet_leaf_34_clk),
    .D(net509),
    .RESET_B(clknet_1_0__leaf_net1160),
    .SCD(net1185),
    .SCE(clknet_1_1__leaf_net1150),
    .SET_B(net1240),
    .Q(net1157),
    .Q_N(net513));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(net512),
    .A1(clknet_1_0__leaf_net1150),
    .A2(clknet_1_0__leaf_net1160),
    .A3(net1185),
    .S0(net1000),
    .S1(net1049),
    .X(net514));
 sky130_fd_sc_hd__mux4_1 c492 (.A0(net512),
    .A1(net347),
    .A2(clknet_1_0__leaf_net1160),
    .A3(net1185),
    .S0(clknet_1_0__leaf_net1150),
    .S1(net1053),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(net1161),
    .A1(clknet_1_0__leaf_net1150),
    .A2(net1185),
    .A3(clknet_1_1__leaf_net1160),
    .S0(net822),
    .S1(net1020),
    .X(net516));
 sky130_fd_sc_hd__sdfbbn_1 c494 (.CLK_N(clknet_leaf_34_clk),
    .D(net510),
    .RESET_B(net1185),
    .SCD(clknet_1_0__leaf_net1160),
    .SCE(clknet_1_1__leaf_net1150),
    .SET_B(net1241),
    .Q(net518),
    .Q_N(net517));
 sky130_fd_sc_hd__a2111o_1 c495 (.A1(net518),
    .A2(net1185),
    .B1(clknet_1_0__leaf_net1150),
    .C1(clknet_1_1__leaf_net1160),
    .D1(net1056),
    .X(net519));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(net518),
    .A1(net1185),
    .A2(clknet_1_0__leaf_net1150),
    .A3(clknet_1_1__leaf_net1160),
    .S0(net1054),
    .S1(net1055),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net1157),
    .A1(net1185),
    .A2(clknet_1_1__leaf_net1160),
    .A3(clknet_1_1__leaf_net1150),
    .S0(net821),
    .S1(net1241),
    .X(net521));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(clknet_1_1__leaf_net1160),
    .A1(clknet_1_0__leaf_net1150),
    .A2(net861),
    .A3(net1020),
    .S0(net1055),
    .S1(net1058),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(net517),
    .A1(net1020),
    .A2(net1054),
    .A3(net1055),
    .S0(net1057),
    .S1(net1059),
    .X(net523));
 sky130_fd_sc_hd__or4bb_1 c50 (.A(net18),
    .B(net25),
    .C_N(net1166),
    .D_N(net1174),
    .X(net26));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(net513),
    .A1(net1185),
    .A2(net1020),
    .A3(clknet_1_0__leaf_net1050),
    .S0(net1057),
    .S1(net1059),
    .X(net524));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(net523),
    .A1(clknet_1_1__leaf_net1160),
    .A2(clknet_1_1__leaf_net524),
    .A3(net1056),
    .S0(net1058),
    .S1(net1059),
    .X(net525));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(net523),
    .A1(clknet_1_0__leaf_net524),
    .A2(clknet_1_1__leaf_net1160),
    .A3(net978),
    .S0(net1059),
    .S1(net1148),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(clknet_1_0__leaf_net524),
    .A1(net523),
    .A2(net1162),
    .A3(net1058),
    .S0(net1059),
    .S1(net1148),
    .X(net1147));
 sky130_fd_sc_hd__and2_2 c504 (.A(net413),
    .B(net1192),
    .X(net527));
 sky130_fd_sc_hd__buf_1 c505 (.A(net766),
    .X(net528));
 sky130_fd_sc_hd__buf_1 c506 (.A(net766),
    .X(net529));
 sky130_fd_sc_hd__clkbuf_1 c507 (.X(net530));
 sky130_fd_sc_hd__and2_0 c508 (.A(net528),
    .B(net1192),
    .X(net531));
 sky130_fd_sc_hd__clkbuf_2 c509 (.A(net795),
    .X(net532));
 sky130_fd_sc_hd__sdfbbn_1 c51 (.CLK_N(clknet_leaf_1_clk),
    .D(net22),
    .RESET_B(net24),
    .SCD(net25),
    .SCE(net1174),
    .SET_B(net21),
    .Q(net28),
    .Q_N(net27));
 sky130_fd_sc_hd__buf_1 c510 (.A(clknet_1_1__leaf_net1128),
    .X(net533));
 sky130_fd_sc_hd__sdfstp_1 c511 (.CLK(clknet_leaf_13_clk),
    .D(net531),
    .SCD(net529),
    .SCE(clknet_1_0__leaf_net533),
    .SET_B(net527),
    .Q(net534));
 sky130_fd_sc_hd__and2_0 c512 (.A(clknet_1_0__leaf_net533),
    .B(net531),
    .X(net535));
 sky130_fd_sc_hd__a2111o_1 c513 (.A1(net529),
    .A2(net534),
    .B1(clknet_1_0__leaf_net535),
    .C1(net1192),
    .D1(net527),
    .X(net536));
 sky130_fd_sc_hd__sdfbbp_1 c514 (.CLK(clknet_leaf_12_clk),
    .D(net1270),
    .RESET_B(net413),
    .SCD(clknet_1_0__leaf_net535),
    .SCE(net527),
    .SET_B(net1226),
    .Q(net538),
    .Q_N(net537));
 sky130_fd_sc_hd__and2_0 c515 (.A(net538),
    .B(clknet_1_1__leaf_net535),
    .X(net539));
 sky130_fd_sc_hd__mux4_1 c516 (.A0(clknet_1_0__leaf_net533),
    .A1(clknet_1_0__leaf_net539),
    .A2(net537),
    .A3(clknet_1_1__leaf_net535),
    .S0(net532),
    .S1(net817),
    .X(net540));
 sky130_fd_sc_hd__mux4_1 c517 (.A0(net532),
    .A1(clknet_1_0__leaf_net535),
    .A2(clknet_1_0__leaf_net539),
    .A3(net537),
    .S0(net1191),
    .S1(net1060),
    .X(net541));
 sky130_fd_sc_hd__mux4_1 c518 (.A0(clknet_1_1__leaf_net535),
    .A1(net538),
    .A2(clknet_1_0__leaf_net539),
    .A3(net527),
    .S0(net1060),
    .S1(net1215),
    .X(net542));
 sky130_fd_sc_hd__mux4_1 c519 (.A0(net527),
    .A1(net537),
    .A2(net532),
    .A3(net817),
    .S0(net1060),
    .S1(net1061),
    .X(net543));
 sky130_fd_sc_hd__mux4_1 c52 (.A0(net23),
    .A1(net28),
    .A2(net1166),
    .A3(net1174),
    .S0(net25),
    .X(net29));
 sky130_fd_sc_hd__mux4_1 c520 (.A0(net529),
    .A1(clknet_1_1__leaf_net539),
    .A2(net534),
    .A3(net527),
    .S0(net1060),
    .S1(net1062),
    .X(net544));
 sky130_fd_sc_hd__mux4_1 c521 (.A0(net532),
    .A1(clknet_1_1__leaf_net539),
    .A2(net817),
    .A3(net1060),
    .S0(net1062),
    .S1(net1064),
    .X(net545));
 sky130_fd_sc_hd__mux4_1 c522 (.A0(net532),
    .A1(net527),
    .A2(net538),
    .A3(net1062),
    .S0(net1063),
    .S1(net1278),
    .X(net546));
 sky130_fd_sc_hd__mux4_1 c523 (.A0(clknet_1_1__leaf_net539),
    .A1(clknet_1_1__leaf_net533),
    .A2(net534),
    .A3(net1062),
    .S0(net1064),
    .S1(net1067),
    .X(net547));
 sky130_fd_sc_hd__mux4_1 c524 (.A0(clknet_1_1__leaf_net533),
    .A1(net1025),
    .A2(net1060),
    .A3(net1063),
    .S0(net1066),
    .S1(net1067),
    .X(net548));
 sky130_fd_sc_hd__and2_0 c525 (.A(clknet_1_0__leaf_net548),
    .B(net825),
    .X(net549));
 sky130_fd_sc_hd__and2_0 c526 (.A(clknet_1_0__leaf_net549),
    .B(net1196),
    .X(net550));
 sky130_fd_sc_hd__buf_1 c527 (.A(net790),
    .X(net551));
 sky130_fd_sc_hd__and2_2 c528 (.A(net551),
    .B(net1068),
    .X(net552));
 sky130_fd_sc_hd__and3_1 c529 (.A(net552),
    .B(net551),
    .C(clknet_1_0__leaf_net548),
    .X(net553));
 sky130_fd_sc_hd__a2111o_1 c53 (.A1(net19),
    .A2(net1166),
    .B1(net25),
    .C1(net1174),
    .D1(net837),
    .X(net30));
 sky130_fd_sc_hd__and3_1 c530 (.A(clknet_1_1__leaf_net549),
    .B(net552),
    .C(clknet_1_0__leaf_net553),
    .X(net554));
 sky130_fd_sc_hd__sdfbbn_1 c531 (.CLK_N(clknet_leaf_14_clk),
    .D(clknet_1_0__leaf_net554),
    .RESET_B(clknet_1_1__leaf_net549),
    .SCD(net552),
    .SCE(clknet_1_0__leaf_net553),
    .SET_B(net1196),
    .Q(net556),
    .Q_N(net555));
 sky130_fd_sc_hd__sdfbbn_1 c532 (.CLK_N(clknet_leaf_14_clk),
    .D(net1249),
    .RESET_B(clknet_1_0__leaf_net548),
    .SCD(clknet_1_0__leaf_net554),
    .SCE(net551),
    .SET_B(net1024),
    .Q(net558),
    .Q_N(net557));
 sky130_fd_sc_hd__sdfbbp_1 c533 (.CLK(clknet_leaf_14_clk),
    .D(net551),
    .RESET_B(net1227),
    .SCD(clknet_1_0__leaf_net553),
    .SCE(clknet_1_0__leaf_net548),
    .SET_B(clknet_1_1__leaf_net554),
    .Q(net560),
    .Q_N(net559));
 sky130_fd_sc_hd__mux4_1 c534 (.A0(net556),
    .A1(clknet_1_0__leaf_net553),
    .A2(net551),
    .A3(clknet_1_0__leaf_net554),
    .S0(net552),
    .S1(net1068),
    .X(net561));
 sky130_fd_sc_hd__sdfbbn_1 c535 (.CLK_N(clknet_leaf_18_clk),
    .D(net1227),
    .RESET_B(clknet_1_1__leaf_net554),
    .SCD(net552),
    .SCE(clknet_1_0__leaf_net553),
    .SET_B(clknet_1_0__leaf_net550),
    .Q(net563),
    .Q_N(net562));
 sky130_fd_sc_hd__mux4_1 c536 (.A0(net552),
    .A1(clknet_1_0__leaf_net554),
    .A2(clknet_1_0__leaf_net553),
    .A3(net562),
    .S0(net555),
    .S1(clknet_1_0__leaf_net549),
    .X(net564));
 sky130_fd_sc_hd__mux4_1 c537 (.A0(net563),
    .A1(net551),
    .A2(clknet_1_1__leaf_net553),
    .A3(clknet_1_1__leaf_net554),
    .S0(net559),
    .S1(net1069),
    .X(net565));
 sky130_fd_sc_hd__sdfbbn_1 c538 (.CLK_N(clknet_leaf_16_clk),
    .D(clknet_1_1__leaf_net554),
    .RESET_B(net562),
    .SCD(clknet_1_0__leaf_net553),
    .SCE(net557),
    .SET_B(clknet_1_0__leaf_net1070),
    .Q(net567),
    .Q_N(net566));
 sky130_fd_sc_hd__mux4_1 c539 (.A0(clknet_1_1__leaf_net553),
    .A1(net563),
    .A2(net552),
    .A3(clknet_1_1__leaf_net554),
    .S0(net818),
    .S1(clknet_1_1__leaf_net1070),
    .X(net568));
 sky130_fd_sc_hd__mux4_1 c54 (.A0(net28),
    .A1(net25),
    .A2(net1166),
    .A3(net1174),
    .S0(net837),
    .S1(net889),
    .X(net31));
 sky130_fd_sc_hd__mux4_1 c540 (.A0(net567),
    .A1(net563),
    .A2(clknet_1_1__leaf_net554),
    .A3(net560),
    .S0(clknet_1_0__leaf_net1070),
    .S1(clknet_1_0__leaf_net1071),
    .X(net569));
 sky130_fd_sc_hd__mux4_1 c541 (.A0(net563),
    .A1(net566),
    .A2(net552),
    .A3(clknet_1_1__leaf_net553),
    .S0(clknet_1_0__leaf_net1071),
    .S1(clknet_1_0__leaf_net1072),
    .X(net570));
 sky130_fd_sc_hd__mux4_1 c542 (.A0(clknet_1_1__leaf_net550),
    .A1(net562),
    .A2(clknet_1_0__leaf_net570),
    .A3(net552),
    .S0(clknet_1_0__leaf_net1071),
    .S1(clknet_1_0__leaf_net1072),
    .X(net571));
 sky130_fd_sc_hd__mux4_1 c543 (.A0(clknet_1_0__leaf_net570),
    .A1(net1069),
    .A2(clknet_1_1__leaf_net1070),
    .A3(clknet_1_1__leaf_net1071),
    .S0(clknet_1_0__leaf_net1072),
    .S1(net1074),
    .X(net572));
 sky130_fd_sc_hd__mux4_1 c544 (.A0(net560),
    .A1(clknet_1_1__leaf_net570),
    .A2(net567),
    .A3(net562),
    .S0(net885),
    .S1(clknet_1_1__leaf_net1072),
    .X(net573));
 sky130_fd_sc_hd__mux4_1 c545 (.A0(clknet_1_1__leaf_net553),
    .A1(net818),
    .A2(net885),
    .A3(clknet_1_1__leaf_net1070),
    .S0(clknet_1_1__leaf_net1071),
    .S1(clknet_1_1__leaf_net1072),
    .X(net574));
 sky130_fd_sc_hd__and2_0 c546 (.A(net1029),
    .B(net1073),
    .X(net575));
 sky130_fd_sc_hd__and2_2 c547 (.A(net1036),
    .B(net1196),
    .X(net576));
 sky130_fd_sc_hd__and2_1 c548 (.A(net436),
    .B(net1198),
    .X(net577));
 sky130_fd_sc_hd__and2_0 c549 (.A(net575),
    .B(net576),
    .X(net578));
 sky130_fd_sc_hd__mux4_1 c55 (.A0(net24),
    .A1(net1174),
    .A2(net25),
    .A3(net27),
    .S0(net1166),
    .S1(net889),
    .X(net32));
 sky130_fd_sc_hd__and3_1 c550 (.A(net1172),
    .B(net1029),
    .C(net1074),
    .X(net579));
 sky130_fd_sc_hd__sdfstp_1 c551 (.CLK(clknet_leaf_17_clk),
    .D(net576),
    .SCD(clknet_1_0__leaf_net574),
    .SCE(net1172),
    .SET_B(net577),
    .Q(net580));
 sky130_fd_sc_hd__and3_1 c552 (.A(net1173),
    .B(net576),
    .C(net1036),
    .X(net581));
 sky130_fd_sc_hd__and3_1 c553 (.A(net577),
    .B(net1173),
    .C(net1036),
    .X(net582));
 sky130_fd_sc_hd__buf_1 c554 (.A(net803),
    .X(net583));
 sky130_fd_sc_hd__mux4_1 c555 (.A0(net579),
    .A1(net580),
    .A2(net583),
    .A3(net1172),
    .S0(net576),
    .S1(net582),
    .X(net584));
 sky130_fd_sc_hd__mux4_2 c556 (.A0(net577),
    .A1(net583),
    .A2(net580),
    .A3(net1172),
    .S0(net576),
    .S1(net1076),
    .X(net585));
 sky130_fd_sc_hd__mux4_1 c557 (.A0(net582),
    .A1(net577),
    .A2(net583),
    .A3(net1172),
    .S0(net585),
    .S1(net1076),
    .X(net586));
 sky130_fd_sc_hd__mux4_1 c558 (.A0(net581),
    .A1(net585),
    .A2(net1173),
    .A3(net580),
    .S0(net1075),
    .S1(net1078),
    .X(net587));
 sky130_fd_sc_hd__mux4_1 c559 (.A0(net306),
    .A1(net585),
    .A2(net1173),
    .A3(net1029),
    .S0(net1076),
    .S1(net1077),
    .X(net588));
 sky130_fd_sc_hd__mux4_1 c56 (.A0(net22),
    .A1(net28),
    .A2(net25),
    .A3(net1166),
    .S0(net20),
    .S1(clknet_1_1__leaf_net904),
    .X(net33));
 sky130_fd_sc_hd__mux4_1 c560 (.A0(net577),
    .A1(net582),
    .A2(net1173),
    .A3(net883),
    .S0(net1075),
    .S1(net1079),
    .X(net589));
 sky130_fd_sc_hd__mux4_1 c561 (.A0(net583),
    .A1(net585),
    .A2(net1172),
    .A3(net1075),
    .S0(net1078),
    .S1(net1080),
    .X(net590));
 sky130_fd_sc_hd__mux4_1 c562 (.A0(net582),
    .A1(net1172),
    .A2(net1076),
    .A3(net1078),
    .S0(net1079),
    .S1(net1080),
    .X(net591));
 sky130_fd_sc_hd__mux4_1 c563 (.A0(net580),
    .A1(net1173),
    .A2(net582),
    .A3(net1076),
    .S0(net1079),
    .S1(net1082),
    .X(net592));
 sky130_fd_sc_hd__mux4_1 c564 (.A0(net576),
    .A1(net585),
    .A2(net883),
    .A3(net1079),
    .S0(net1080),
    .S1(net1082),
    .X(net593));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net585),
    .A1(clknet_1_1__leaf_net891),
    .A2(net1075),
    .A3(net1080),
    .S0(net1081),
    .S1(net1082),
    .X(net594));
 sky130_fd_sc_hd__mux4_2 c566 (.A0(net859),
    .A1(clknet_1_1__leaf_net891),
    .A2(net1077),
    .A3(net1079),
    .S0(net1080),
    .S1(net1082),
    .X(net595));
 sky130_fd_sc_hd__a2111o_1 c567 (.A1(net576),
    .A2(clknet_1_0__leaf_net595),
    .B1(net1173),
    .C1(net1197),
    .D1(net1196),
    .X(net596));
 sky130_fd_sc_hd__buf_1 c568 (.A(net885),
    .X(net597));
 sky130_fd_sc_hd__sdfbbp_1 c569 (.CLK(clknet_leaf_28_clk),
    .D(net597),
    .RESET_B(clknet_1_0__leaf_net596),
    .SCD(net1197),
    .SCE(net1081),
    .SET_B(net1082),
    .Q(net599),
    .Q_N(net598));
 sky130_fd_sc_hd__mux4_1 c57 (.A0(net28),
    .A1(net25),
    .A2(net1166),
    .A3(net1174),
    .S0(clknet_1_0__leaf_net904),
    .S1(clknet_1_0__leaf_net906),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 c570 (.A(net885),
    .X(net600));
 sky130_fd_sc_hd__sdfbbn_1 c571 (.CLK_N(clknet_leaf_29_clk),
    .D(net597),
    .RESET_B(net599),
    .SCD(clknet_1_0__leaf_net596),
    .SCE(net600),
    .SET_B(net1259),
    .Q(net602),
    .Q_N(net601));
 sky130_fd_sc_hd__mux4_1 c572 (.A0(net576),
    .A1(net600),
    .A2(net598),
    .A3(net601),
    .S0(clknet_1_0__leaf_net596),
    .S1(net1196),
    .X(net603));
 sky130_fd_sc_hd__mux4_1 c573 (.A0(net599),
    .A1(net602),
    .A2(net600),
    .A3(net597),
    .S0(net1036),
    .S1(net1083),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 c574 (.A0(net597),
    .A1(net600),
    .A2(clknet_1_0__leaf_net596),
    .A3(net1197),
    .S0(net1081),
    .S1(net1083),
    .X(net605));
 sky130_fd_sc_hd__mux4_1 c575 (.A0(clknet_1_0__leaf_net596),
    .A1(net602),
    .A2(net598),
    .A3(net1197),
    .S0(net1083),
    .S1(net1085),
    .X(net606));
 sky130_fd_sc_hd__mux4_1 c576 (.A0(net325),
    .A1(net1173),
    .A2(net601),
    .A3(clknet_1_1__leaf_net596),
    .S0(net1083),
    .S1(net1087),
    .X(net607));
 sky130_fd_sc_hd__mux4_1 c577 (.A0(net597),
    .A1(net601),
    .A2(clknet_1_0__leaf_net848),
    .A3(net1083),
    .S0(net1085),
    .S1(net1087),
    .X(net608));
 sky130_fd_sc_hd__mux4_1 c578 (.A0(net600),
    .A1(clknet_1_0__leaf_net608),
    .A2(clknet_1_1__leaf_net596),
    .A3(clknet_1_0__leaf_net848),
    .S0(net1084),
    .S1(net1087),
    .X(net609));
 sky130_fd_sc_hd__mux4_1 c579 (.A0(net602),
    .A1(clknet_1_0__leaf_net608),
    .A2(net599),
    .A3(clknet_1_1__leaf_net596),
    .S0(net1087),
    .S1(net1088),
    .X(net610));
 sky130_fd_sc_hd__mux4_1 c58 (.A0(net27),
    .A1(net25),
    .A2(net837),
    .A3(clknet_1_0__leaf_net904),
    .S0(clknet_1_1__leaf_net906),
    .S1(net908),
    .X(net35));
 sky130_fd_sc_hd__mux4_1 c580 (.A0(net323),
    .A1(net600),
    .A2(clknet_1_1__leaf_net596),
    .A3(clknet_1_1__leaf_net892),
    .S0(net1083),
    .S1(net1088),
    .X(net611));
 sky130_fd_sc_hd__mux4_2 c581 (.A0(net604),
    .A1(net601),
    .A2(net1084),
    .A3(net1086),
    .S0(net1088),
    .S1(net1089),
    .X(net612));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(net612),
    .A1(clknet_1_1__leaf_net892),
    .A2(net1082),
    .A3(net1084),
    .S0(net1088),
    .S1(net1089),
    .X(net1153));
 sky130_fd_sc_hd__mux4_1 c583 (.A0(net600),
    .A1(net612),
    .A2(clknet_1_0__leaf_net1153),
    .A3(clknet_1_1__leaf_net608),
    .S0(net1088),
    .S1(net1089),
    .X(net613));
 sky130_fd_sc_hd__mux4_1 c584 (.A0(clknet_1_1__leaf_net608),
    .A1(clknet_1_0__leaf_net1153),
    .A2(net599),
    .A3(net1086),
    .S0(net1088),
    .S1(net1089),
    .X(net614));
 sky130_fd_sc_hd__mux4_1 c585 (.A0(clknet_1_1__leaf_net608),
    .A1(net1085),
    .A2(net1088),
    .A3(net1089),
    .S0(net1090),
    .S1(clknet_1_0__leaf_net1091),
    .X(net615));
 sky130_fd_sc_hd__mux4_1 c586 (.A0(clknet_1_1__leaf_net615),
    .A1(net1197),
    .A2(net1085),
    .A3(net1086),
    .S0(net1090),
    .S1(clknet_1_0__leaf_net1091),
    .X(net616));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(net616),
    .A1(clknet_1_0__leaf_net1153),
    .A2(net602),
    .A3(clknet_1_0__leaf_net615),
    .S0(net1089),
    .S1(clknet_1_1__leaf_net1091),
    .X(net617));
 sky130_fd_sc_hd__and2_4 c588 (.A(clknet_1_1__leaf_net595),
    .B(net1090),
    .X(net618));
 sky130_fd_sc_hd__and2_4 c589 (.A(clknet_1_0__leaf_net618),
    .B(net1156),
    .X(net619));
 sky130_fd_sc_hd__mux4_1 c59 (.A0(net25),
    .A1(clknet_1_0__leaf_net35),
    .A2(net28),
    .A3(net1166),
    .S0(clknet_1_0__leaf_net906),
    .S1(net907),
    .X(net36));
 sky130_fd_sc_hd__buf_1 c590 (.A(net875),
    .X(net620));
 sky130_fd_sc_hd__dlymetal6s2s_1 c591 (.A(net875),
    .X(net621));
 sky130_fd_sc_hd__or4bb_1 c592 (.A(net621),
    .B(net1212),
    .C_N(net1184),
    .D_N(clknet_1_0__leaf_net619),
    .X(net622));
 sky130_fd_sc_hd__sdfbbn_1 c593 (.CLK_N(clknet_leaf_26_clk),
    .D(net621),
    .RESET_B(net1269),
    .SCD(clknet_1_1__leaf_net619),
    .SCE(clknet_1_1__leaf_net618),
    .SET_B(net1090),
    .Q(net624),
    .Q_N(net623));
 sky130_fd_sc_hd__mux4_1 c594 (.A0(clknet_1_0__leaf_net619),
    .A1(net623),
    .A2(net1184),
    .A3(net1212),
    .S0(net621),
    .S1(net827),
    .X(net625));
 sky130_fd_sc_hd__sdfbbp_1 c595 (.CLK(clknet_leaf_26_clk),
    .D(net1184),
    .RESET_B(clknet_1_1__leaf_net618),
    .SCD(clknet_1_1__leaf_net619),
    .SCE(net623),
    .SET_B(net883),
    .Q(net627),
    .Q_N(net626));
 sky130_fd_sc_hd__mux4_1 c596 (.A0(clknet_1_0__leaf_net619),
    .A1(clknet_1_0__leaf_net618),
    .A2(net1184),
    .A3(net626),
    .S0(net828),
    .S1(clknet_1_1__leaf_net1050),
    .X(net628));
 sky130_fd_sc_hd__mux4_1 c597 (.A0(net612),
    .A1(net624),
    .A2(clknet_1_0__leaf_net618),
    .A3(net626),
    .S0(net1184),
    .S1(clknet_1_0__leaf_net619),
    .X(net629));
 sky130_fd_sc_hd__mux4_1 c598 (.A0(net1184),
    .A1(net627),
    .A2(clknet_1_0__leaf_net619),
    .A3(net621),
    .S0(net1212),
    .S1(clknet_1_0__leaf_net1092),
    .X(net630));
 sky130_fd_sc_hd__mux4_2 c599 (.A0(net1184),
    .A1(net621),
    .A2(clknet_1_0__leaf_net618),
    .A3(clknet_1_0__leaf_net619),
    .S1(clknet_1_0__leaf_net1092),
    .X(net886));
 sky130_fd_sc_hd__mux4_1 c60 (.A0(clknet_1_1__leaf_net35),
    .A1(net24),
    .A2(net27),
    .A3(clknet_1_1__leaf_net906),
    .S0(net908),
    .S1(net910),
    .X(net37));
 sky130_fd_sc_hd__mux4_1 c600 (.A0(net627),
    .A1(net621),
    .A2(net620),
    .A3(clknet_1_1__leaf_net619),
    .S0(clknet_1_0__leaf_net886),
    .S1(clknet_1_1__leaf_net1092),
    .X(net632));
 sky130_fd_sc_hd__mux4_1 c601 (.A0(net627),
    .A1(net621),
    .A2(net623),
    .A3(net1184),
    .S0(clknet_1_0__leaf_net618),
    .S1(clknet_1_0__leaf_net1092),
    .X(net633));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(net624),
    .A1(net627),
    .A2(clknet_1_1__leaf_net1153),
    .A3(clknet_1_1__leaf_net618),
    .S0(net878),
    .S1(clknet_1_1__leaf_net1092),
    .X(net634));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(net624),
    .A1(net633),
    .A2(clknet_1_1__leaf_net618),
    .A3(net1184),
    .S0(clknet_1_1__leaf_net1092),
    .S1(clknet_1_0__leaf_net1093),
    .X(net635));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(net620),
    .A1(net1212),
    .A2(net828),
    .A3(clknet_1_0__leaf_net1092),
    .S0(clknet_1_0__leaf_net1093),
    .S1(net1094),
    .X(net636));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(clknet_1_1__leaf_net618),
    .A1(clknet_1_1__leaf_net619),
    .A2(net864),
    .A3(clknet_1_1__leaf_net1092),
    .S0(clknet_1_1__leaf_net1093),
    .S1(net1155),
    .X(net637));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net636),
    .A1(clknet_1_1__leaf_net619),
    .A2(net864),
    .A3(net883),
    .S0(clknet_1_1__leaf_net886),
    .S1(net1095),
    .X(net638));
 sky130_fd_sc_hd__mux4_2 c607 (.A0(net624),
    .A1(net874),
    .A2(net878),
    .A3(clknet_1_0__leaf_net886),
    .S0(clknet_1_1__leaf_net1093),
    .S1(net1096),
    .X(net639));
 sky130_fd_sc_hd__mux4_2 c608 (.A0(net639),
    .A1(net626),
    .A2(net612),
    .A3(net874),
    .S0(clknet_1_1__leaf_net1093),
    .S1(net1096),
    .X(net1154));
 sky130_fd_sc_hd__mux4_1 c61 (.A0(net19),
    .A1(clknet_1_0__leaf_net35),
    .A2(clknet_1_0__leaf_net37),
    .A3(net27),
    .S0(clknet_1_1__leaf_net906),
    .S1(net909),
    .X(net38));
 sky130_fd_sc_hd__mux4_1 c62 (.A0(clknet_1_1__leaf_net37),
    .A1(net38),
    .A2(clknet_1_1__leaf_net35),
    .A3(net21),
    .S0(net908),
    .S1(net910),
    .X(net39));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(clknet_1_0__leaf_net1154),
    .A1(clknet_1_1__leaf_net1150),
    .A2(net1162),
    .A3(clknet_1_1__leaf_net848),
    .S0(net978),
    .S1(net1240),
    .X(net640));
 sky130_fd_sc_hd__and2_0 c63 (.A(net1180),
    .B(net43),
    .X(net40));
 sky130_fd_sc_hd__and2_0 c630 (.A(clknet_1_1__leaf_net548),
    .B(net1196),
    .X(net641));
 sky130_fd_sc_hd__and2_0 c631 (.A(clknet_1_0__leaf_net641),
    .B(net1025),
    .X(net642));
 sky130_fd_sc_hd__clkbuf_1 c632 (.A(net872),
    .X(net643));
 sky130_fd_sc_hd__buf_1 c633 (.A(net872),
    .X(net644));
 sky130_fd_sc_hd__sedfxbp_1 c634 (.CLK(clknet_leaf_13_clk),
    .D(net1182),
    .DE(clknet_1_0__leaf_net548),
    .SCD(clknet_1_0__leaf_net642),
    .SCE(net1181),
    .Q(net646),
    .Q_N(net645));
 sky130_fd_sc_hd__sedfxbp_1 c635 (.CLK(clknet_leaf_18_clk),
    .D(net1272),
    .DE(clknet_1_0__leaf_net642),
    .SCD(net1181),
    .SCE(net1182),
    .Q(net648),
    .Q_N(net647));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(clknet_1_0__leaf_net641),
    .A1(net647),
    .A2(net1181),
    .A3(net1182),
    .S0(clknet_1_0__leaf_net642),
    .S1(net1023),
    .X(net649));
 sky130_fd_sc_hd__sdfbbn_1 c637 (.CLK_N(clknet_leaf_18_clk),
    .D(net648),
    .RESET_B(net1182),
    .SCD(clknet_1_0__leaf_net642),
    .SCE(net1181),
    .SET_B(net1234),
    .Q(net651),
    .Q_N(net650));
 sky130_fd_sc_hd__sdfbbn_1 c638 (.CLK_N(clknet_leaf_18_clk),
    .D(net1252),
    .RESET_B(clknet_1_1__leaf_net641),
    .SCD(clknet_1_0__leaf_net642),
    .SCE(net1181),
    .SET_B(net1183),
    .Q(net653),
    .Q_N(net652));
 sky130_fd_sc_hd__a2111o_1 c639 (.A1(net653),
    .A2(net650),
    .B1(clknet_1_0__leaf_net642),
    .C1(net1181),
    .D1(net1182),
    .X(net654));
 sky130_fd_sc_hd__and2_1 c64 (.A(net43),
    .B(net1180),
    .X(net41));
 sky130_fd_sc_hd__sdfbbp_1 c640 (.CLK(clknet_leaf_18_clk),
    .D(clknet_1_0__leaf_net642),
    .RESET_B(net653),
    .SCD(net1181),
    .SCE(net1182),
    .SET_B(net1097),
    .Q(net656),
    .Q_N(net655));
 sky130_fd_sc_hd__mux4_1 c641 (.A0(net645),
    .A1(net1181),
    .A2(net652),
    .A3(clknet_1_0__leaf_net642),
    .S0(net1182),
    .S1(net1097),
    .X(net657));
 sky130_fd_sc_hd__mux4_1 c642 (.A0(net653),
    .A1(net655),
    .A2(net1181),
    .A3(net1182),
    .S0(clknet_1_1__leaf_net642),
    .S1(net1205),
    .X(net658));
 sky130_fd_sc_hd__mux4_1 c643 (.A0(net646),
    .A1(net652),
    .A2(clknet_1_1__leaf_net642),
    .A3(net1182),
    .S0(net1205),
    .S1(net1099),
    .X(net659));
 sky130_fd_sc_hd__mux4_1 c644 (.A0(net656),
    .A1(net653),
    .A2(clknet_1_1__leaf_net642),
    .A3(net1181),
    .S0(net1205),
    .S1(net1100),
    .X(net660));
 sky130_fd_sc_hd__mux4_1 c645 (.A0(net648),
    .A1(clknet_1_1__leaf_net642),
    .A2(net652),
    .A3(net877),
    .S0(net1205),
    .S1(net1100),
    .X(net661));
 sky130_fd_sc_hd__mux4_1 c646 (.A0(net651),
    .A1(net655),
    .A2(net653),
    .A3(net1205),
    .S0(net1100),
    .S1(net1101),
    .X(net662));
 sky130_fd_sc_hd__mux4_1 c647 (.A0(net662),
    .A1(net652),
    .A2(net877),
    .A3(net1205),
    .S0(net1099),
    .S1(net1101),
    .X(net663));
 sky130_fd_sc_hd__mux4_1 c648 (.A0(net644),
    .A1(net656),
    .A2(net662),
    .A3(net663),
    .S0(net1196),
    .S1(net1101),
    .X(net664));
 sky130_fd_sc_hd__mux4_1 c649 (.A0(net663),
    .A1(net662),
    .A2(net1183),
    .A3(net644),
    .S0(net1099),
    .S1(net1101),
    .X(net665));
 sky130_fd_sc_hd__and2_1 c65 (.A(net1130),
    .B(net1203),
    .X(net42));
 sky130_fd_sc_hd__mux4_1 c650 (.A0(net662),
    .A1(net665),
    .A2(net663),
    .A3(net644),
    .S0(clknet_1_1__leaf_net642),
    .S1(net1101),
    .X(net666));
 sky130_fd_sc_hd__and2_0 c651 (.A(clknet_1_1__leaf_net548),
    .B(net1101),
    .X(net667));
 sky130_fd_sc_hd__and2_0 c652 (.A(net1183),
    .B(clknet_1_0__leaf_net667),
    .X(net668));
 sky130_fd_sc_hd__sedfxtp_1 c653 (.CLK(clknet_leaf_21_clk),
    .D(clknet_1_0__leaf_net668),
    .DE(clknet_1_1__leaf_net574),
    .SCD(clknet_1_0__leaf_net667),
    .SCE(net1205),
    .Q(net669));
 sky130_fd_sc_hd__sdfbbn_1 c654 (.CLK_N(clknet_leaf_21_clk),
    .D(net669),
    .RESET_B(clknet_1_0__leaf_net668),
    .SCD(net1183),
    .SCE(clknet_1_0__leaf_net667),
    .SET_B(net1205),
    .Q(net671),
    .Q_N(net670));
 sky130_fd_sc_hd__sdfbbn_1 c655 (.CLK_N(clknet_leaf_19_clk),
    .D(net670),
    .RESET_B(clknet_1_0__leaf_net667),
    .SCD(clknet_1_0__leaf_net668),
    .SCE(net1098),
    .SET_B(net1101),
    .Q(net673),
    .Q_N(net672));
 sky130_fd_sc_hd__mux4_1 c656 (.A0(net671),
    .A1(net673),
    .A2(clknet_1_0__leaf_net668),
    .A3(net1183),
    .S0(clknet_1_0__leaf_net667),
    .S1(net818),
    .X(net674));
 sky130_fd_sc_hd__mux4_1 c657 (.A0(net664),
    .A1(net669),
    .A2(net670),
    .A3(clknet_1_0__leaf_net668),
    .S0(net1205),
    .S1(net1102),
    .X(net675));
 sky130_fd_sc_hd__mux4_1 c658 (.A0(clknet_1_0__leaf_net667),
    .A1(net673),
    .A2(clknet_1_1__leaf_net668),
    .A3(net1183),
    .S0(net882),
    .S1(net1205),
    .X(net676));
 sky130_fd_sc_hd__mux4_1 c659 (.A0(net399),
    .A1(net672),
    .A2(clknet_1_1__leaf_net668),
    .A3(net1098),
    .S0(net1102),
    .S1(net1105),
    .X(net677));
 sky130_fd_sc_hd__and2_2 c66 (.A(net1180),
    .B(net907),
    .X(net43));
 sky130_fd_sc_hd__mux4_1 c660 (.A0(net673),
    .A1(clknet_1_1__leaf_net668),
    .A2(clknet_1_1__leaf_net667),
    .A3(net670),
    .S0(net888),
    .S1(net1103),
    .X(net678));
 sky130_fd_sc_hd__mux4_1 c661 (.A0(clknet_1_1__leaf_net668),
    .A1(net672),
    .A2(clknet_1_1__leaf_net667),
    .A3(net882),
    .S0(net1103),
    .S1(net1106),
    .X(net679));
 sky130_fd_sc_hd__mux4_1 c662 (.A0(net673),
    .A1(clknet_1_1__leaf_net667),
    .A2(clknet_1_1__leaf_net668),
    .A3(net888),
    .S0(net1102),
    .S1(net1106),
    .X(net680));
 sky130_fd_sc_hd__mux4_1 c663 (.A0(net672),
    .A1(clknet_1_1__leaf_net667),
    .A2(net1183),
    .A3(net882),
    .S0(net1103),
    .S1(net1107),
    .X(net681));
 sky130_fd_sc_hd__mux4_1 c664 (.A0(clknet_1_0__leaf_net667),
    .A1(net669),
    .A2(clknet_1_0__leaf_net668),
    .A3(net673),
    .S0(clknet_1_0__leaf_net681),
    .S1(net872),
    .X(net682));
 sky130_fd_sc_hd__mux4_1 c665 (.A0(clknet_1_1__leaf_net681),
    .A1(clknet_1_1__leaf_net667),
    .A2(clknet_1_1__leaf_net668),
    .A3(net1105),
    .S0(net1106),
    .S1(net1107),
    .X(net683));
 sky130_fd_sc_hd__mux4_1 c666 (.A0(net671),
    .A1(clknet_1_1__leaf_net574),
    .A2(clknet_1_1__leaf_net667),
    .A3(net1104),
    .S0(net1107),
    .S1(net1108),
    .X(net684));
 sky130_fd_sc_hd__mux4_1 c667 (.A0(net671),
    .A1(clknet_1_0__leaf_net681),
    .A2(clknet_1_1__leaf_net668),
    .A3(net1183),
    .S0(net1107),
    .S1(net1108),
    .X(net685));
 sky130_fd_sc_hd__mux4_1 c668 (.A0(clknet_1_1__leaf_net681),
    .A1(net672),
    .A2(net1107),
    .A3(net1108),
    .S0(clknet_1_0__leaf_net1109),
    .S1(clknet_1_1__leaf_net1110),
    .X(net686));
 sky130_fd_sc_hd__mux4_1 c669 (.A0(clknet_1_1__leaf_net667),
    .A1(clknet_1_0__leaf_net681),
    .A2(net872),
    .A3(clknet_1_0__leaf_net1109),
    .S0(clknet_1_0__leaf_net1110),
    .S1(clknet_1_0__leaf_net1111),
    .X(net687));
 sky130_fd_sc_hd__dlymetal6s2s_1 c67 (.A(net1126),
    .X(net44));
 sky130_fd_sc_hd__mux4_1 c670 (.A0(clknet_1_1__leaf_net681),
    .A1(net1104),
    .A2(net1107),
    .A3(clknet_1_1__leaf_net1109),
    .S0(clknet_1_1__leaf_net1110),
    .S1(clknet_1_1__leaf_net1111),
    .X(net688));
 sky130_fd_sc_hd__mux4_1 c671 (.A0(net669),
    .A1(net869),
    .A2(net882),
    .A3(net1107),
    .S0(clknet_1_0__leaf_net1110),
    .S1(clknet_1_0__leaf_net1111),
    .X(net689));
 sky130_fd_sc_hd__and2_1 c672 (.A(net1172),
    .B(net1080),
    .X(net690));
 sky130_fd_sc_hd__buf_1 c673 (.A(net775),
    .X(net691));
 sky130_fd_sc_hd__and2_0 c674 (.A(net691),
    .B(net1214),
    .X(net692));
 sky130_fd_sc_hd__clkbuf_1 c675 (.A(net775),
    .X(net693));
 sky130_fd_sc_hd__and2_0 c676 (.A(clknet_1_0__leaf_net692),
    .B(net691),
    .X(net694));
 sky130_fd_sc_hd__and2_1 c677 (.A(net693),
    .B(net691),
    .X(net695));
 sky130_fd_sc_hd__buf_1 c678 (.A(net804),
    .X(net696));
 sky130_fd_sc_hd__buf_1 c679 (.X(net806));
 sky130_fd_sc_hd__and2_0 c68 (.A(net44),
    .B(net1180),
    .X(net45));
 sky130_fd_sc_hd__sdfbbp_1 c680 (.CLK(clknet_leaf_17_clk),
    .D(net690),
    .RESET_B(clknet_1_1__leaf_net694),
    .SCD(net693),
    .SCE(clknet_1_1__leaf_net692),
    .SET_B(net695),
    .Q(net699),
    .Q_N(net698));
 sky130_fd_sc_hd__and2_0 c681 (.A(net691),
    .B(net695),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_1 c682 (.A(net876),
    .X(net701));
 sky130_fd_sc_hd__clkbuf_1 c683 (.A(net876),
    .X(net702));
 sky130_fd_sc_hd__buf_1 c684 (.A(net805),
    .X(net703));
 sky130_fd_sc_hd__mux4_1 c685 (.A0(net701),
    .A1(net690),
    .A2(net703),
    .A3(net1172),
    .S0(net696),
    .S1(clknet_1_1__leaf_net689),
    .X(net704));
 sky130_fd_sc_hd__and3_1 c686 (.A(net703),
    .B(net1080),
    .C(net1081),
    .X(net705));
 sky130_fd_sc_hd__sedfxtp_1 c687 (.CLK(clknet_leaf_21_clk),
    .D(net697),
    .DE(net690),
    .SCD(net696),
    .SCE(clknet_1_1__leaf_net694),
    .Q(net706));
 sky130_fd_sc_hd__and3_1 c688 (.A(net706),
    .B(net697),
    .C(net699),
    .X(net707));
 sky130_fd_sc_hd__or4bb_1 c689 (.A(net707),
    .B(net706),
    .C_N(net695),
    .D_N(clknet_1_1__leaf_net694),
    .X(net708));
 sky130_fd_sc_hd__and3_2 c69 (.A(net42),
    .B(net45),
    .C(net1203),
    .X(net46));
 sky130_fd_sc_hd__mux4_1 c690 (.A0(net705),
    .A1(net703),
    .A2(net706),
    .A3(clknet_1_0__leaf_net694),
    .S0(net819),
    .S1(net1035),
    .X(net709));
 sky130_fd_sc_hd__and3_1 c691 (.A(net706),
    .B(net703),
    .C(net896),
    .X(net710));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(net710),
    .A1(net696),
    .A2(net703),
    .A3(net706),
    .S0(net896),
    .S1(net1082),
    .X(net711));
 sky130_fd_sc_hd__and2_2 c693 (.A(net700),
    .B(net1231),
    .X(net712));
 sky130_fd_sc_hd__buf_2 c694 (.X(net713));
 sky130_fd_sc_hd__clkbuf_2 c695 (.A(net769),
    .X(net714));
 sky130_fd_sc_hd__clkbuf_2 c696 (.X(net715));
 sky130_fd_sc_hd__or4bb_1 c697 (.A(net699),
    .B(clknet_1_0__leaf_net1153),
    .C_N(net1173),
    .D_N(net820),
    .X(net716));
 sky130_fd_sc_hd__clkbuf_1 c698 (.A(net791),
    .X(net717));
 sky130_fd_sc_hd__and3_2 c699 (.A(net717),
    .B(net713),
    .C(net612),
    .X(net718));
 sky130_fd_sc_hd__sdfbbp_1 c70 (.CLK(clknet_leaf_48_clk),
    .D(net40),
    .RESET_B(net44),
    .SCD(net1180),
    .SCE(net43),
    .SET_B(net41),
    .Q(net48),
    .Q_N(net47));
 sky130_fd_sc_hd__sdfbbn_1 c700 (.CLK_N(clknet_leaf_27_clk),
    .D(net712),
    .RESET_B(net715),
    .SCD(net718),
    .SCE(net714),
    .SET_B(net713),
    .Q(net720),
    .Q_N(net719));
 sky130_fd_sc_hd__sdfbbn_1 c701 (.CLK_N(clknet_leaf_27_clk),
    .D(net718),
    .RESET_B(net713),
    .SCD(net1276),
    .SCE(net712),
    .SET_B(net715),
    .Q(net722),
    .Q_N(net721));
 sky130_fd_sc_hd__sdfbbp_1 c702 (.CLK(clknet_leaf_24_clk),
    .D(net702),
    .RESET_B(net718),
    .SCD(net1221),
    .SCE(net714),
    .SET_B(net1228),
    .Q(net724),
    .Q_N(net723));
 sky130_fd_sc_hd__and3_2 c703 (.A(net711),
    .B(net719),
    .C(net714),
    .X(net725));
 sky130_fd_sc_hd__clkbuf_1 c704 (.A(net1120),
    .X(net726));
 sky130_fd_sc_hd__a2111o_1 c705 (.A1(net724),
    .A2(net714),
    .B1(net718),
    .C1(net725),
    .D1(net712),
    .X(net727));
 sky130_fd_sc_hd__or4bb_1 c706 (.A(net1222),
    .B(net725),
    .C_N(net1221),
    .D_N(net718),
    .X(net728));
 sky130_fd_sc_hd__sdfbbn_1 c707 (.CLK_N(clknet_leaf_27_clk),
    .D(net715),
    .RESET_B(net718),
    .SCD(net726),
    .SCE(net712),
    .SET_B(net858),
    .Q(net730),
    .Q_N(net729));
 sky130_fd_sc_hd__sedfxtp_1 c708 (.CLK(clknet_leaf_27_clk),
    .D(net720),
    .DE(net725),
    .SCD(net1228),
    .SCE(net729),
    .Q(net731));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(net720),
    .A1(net714),
    .A2(net1206),
    .A3(net712),
    .S0(net713),
    .S1(net887),
    .X(net732));
 sky130_fd_sc_hd__mux4_1 c71 (.A0(net43),
    .A1(net45),
    .A2(net47),
    .A3(net1180),
    .S0(net46),
    .S1(net907),
    .X(net49));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net725),
    .A1(net1206),
    .A2(net718),
    .A3(net713),
    .S0(net887),
    .S1(net1112),
    .X(net733));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net1228),
    .A1(net1206),
    .A2(net730),
    .A3(net1232),
    .S0(net725),
    .S1(net1113),
    .X(net734));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net731),
    .A1(net725),
    .A2(net718),
    .A3(net870),
    .S0(net895),
    .S1(net1112),
    .X(net735));
 sky130_fd_sc_hd__sdfbbn_1 c713 (.CLK_N(clknet_leaf_23_clk),
    .D(net725),
    .RESET_B(net1206),
    .SCD(net713),
    .SCE(net1113),
    .SET_B(net1233),
    .Q(net737),
    .Q_N(net736));
 sky130_fd_sc_hd__and2_1 c714 (.A(net737),
    .B(net1206),
    .X(net738));
 sky130_fd_sc_hd__buf_1 c715 (.X(net739));
 sky130_fd_sc_hd__and3_1 c716 (.A(net738),
    .B(net736),
    .C(net1206),
    .X(net740));
 sky130_fd_sc_hd__a2111o_1 c717 (.A1(net1219),
    .A2(net612),
    .B1(net738),
    .C1(net1283),
    .D1(net721),
    .X(net741));
 sky130_fd_sc_hd__clkbuf_1 c718 (.A(net777),
    .X(net742));
 sky130_fd_sc_hd__or4bb_4 c719 (.A(net738),
    .B(net1209),
    .C_N(net739),
    .D_N(net820),
    .X(net743));
 sky130_fd_sc_hd__or4bb_1 c72 (.A(net48),
    .B(net43),
    .C_N(net1180),
    .D_N(net44),
    .X(net50));
 sky130_fd_sc_hd__or4bb_1 c720 (.A(net1206),
    .B(net1209),
    .C_N(net743),
    .D_N(net739),
    .X(net744));
 sky130_fd_sc_hd__sdfbbp_1 c721 (.CLK(clknet_leaf_24_clk),
    .D(net730),
    .RESET_B(net743),
    .SCD(net744),
    .SCE(net1206),
    .SET_B(net1209),
    .Q(net746),
    .Q_N(net745));
 sky130_fd_sc_hd__sdfbbn_1 c722 (.CLK_N(clknet_leaf_24_clk),
    .D(net1255),
    .RESET_B(net743),
    .SCD(net744),
    .SCE(net1209),
    .SET_B(net745),
    .Q(net748),
    .Q_N(net747));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net746),
    .A1(net748),
    .A2(net738),
    .A3(net743),
    .S0(net1209),
    .S1(net1090),
    .X(net749));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net748),
    .A1(net1206),
    .A2(net749),
    .A3(net743),
    .S0(net1209),
    .S1(net745),
    .X(net750));
 sky130_fd_sc_hd__a2111o_1 c725 (.A1(net1209),
    .A2(net743),
    .B1(net747),
    .C1(net739),
    .D1(net1117),
    .X(net751));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net751),
    .A1(net748),
    .A2(net740),
    .A3(net743),
    .S0(net1209),
    .S1(net1116),
    .X(net752));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net743),
    .A1(net749),
    .A2(net748),
    .A3(net740),
    .S0(net1209),
    .S1(net1117),
    .X(net753));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net746),
    .A1(net749),
    .A2(net747),
    .S0(net1116),
    .S1(net1118),
    .X(net845));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(net740),
    .A1(net751),
    .A2(net747),
    .A3(net1209),
    .S0(net743),
    .S1(net1117),
    .X(net755));
 sky130_fd_sc_hd__mux4_1 c73 (.A0(net40),
    .A1(net1180),
    .A2(net46),
    .A3(net44),
    .S0(net43),
    .S1(net842),
    .X(net51));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net742),
    .A1(net751),
    .A2(net749),
    .A3(net1116),
    .S0(net1118),
    .S1(net1119),
    .X(net756));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net744),
    .A1(net740),
    .A2(net748),
    .A3(net845),
    .S0(net1119),
    .S1(net1159),
    .X(net757));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(net747),
    .A1(net743),
    .A2(net864),
    .A3(net1116),
    .S0(net1119),
    .S1(net1159),
    .X(net758));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net744),
    .A1(net1115),
    .A2(net1284),
    .A3(net1118),
    .S0(net1119),
    .S1(net1159),
    .X(net759));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(net758),
    .A1(net612),
    .A2(net895),
    .A3(net1117),
    .S0(net1118),
    .S1(net1119),
    .X(net760));
 sky130_fd_sc_hd__mux4_1 c74 (.A0(net41),
    .A1(net50),
    .A2(net43),
    .A3(net42),
    .S0(net907),
    .S1(net912),
    .X(net52));
 sky130_fd_sc_hd__mux4_1 c75 (.A0(net50),
    .A1(net46),
    .A2(net48),
    .A3(net42),
    .S0(net908),
    .S1(net913),
    .X(net53));
 sky130_fd_sc_hd__mux4_1 c76 (.A0(net47),
    .A1(net43),
    .A2(net42),
    .A3(net889),
    .S0(net912),
    .S1(net913),
    .X(net54));
 sky130_fd_sc_hd__mux4_1 c77 (.A0(net45),
    .A1(net48),
    .A2(net54),
    .A3(net1180),
    .S0(net911),
    .S1(net913),
    .X(net55));
 sky130_fd_sc_hd__mux4_1 c78 (.A0(net54),
    .A1(net50),
    .A2(net43),
    .A3(net911),
    .S0(net913),
    .S1(net914),
    .X(net56));
 sky130_fd_sc_hd__mux4_1 c79 (.A0(net44),
    .A1(net46),
    .A2(net911),
    .A3(net913),
    .S0(net914),
    .S1(net915),
    .X(net57));
 sky130_fd_sc_hd__mux4_1 c80 (.A0(net842),
    .A1(net907),
    .A2(net912),
    .A3(net914),
    .S0(net915),
    .S1(net916),
    .X(net58));
 sky130_fd_sc_hd__mux4_2 c81 (.A0(net58),
    .A1(net44),
    .A2(net912),
    .A3(net914),
    .S0(net915),
    .S1(net916),
    .X(net59));
 sky130_fd_sc_hd__mux4_2 c82 (.A0(net59),
    .A1(net58),
    .A2(net47),
    .A3(net44),
    .S0(net915),
    .S1(net916),
    .X(net60));
 sky130_fd_sc_hd__mux4_1 c83 (.A0(net60),
    .A1(net59),
    .A2(net46),
    .A3(net889),
    .S0(net914),
    .S1(net916),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 c84 (.A(net771),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 c85 (.A(net771),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 c86 (.A(net866),
    .X(net64));
 sky130_fd_sc_hd__and2_1 c87 (.A(net1170),
    .B(net64),
    .X(net65));
 sky130_fd_sc_hd__and3_1 c88 (.A(net64),
    .B(net1169),
    .C(net1203),
    .X(net66));
 sky130_fd_sc_hd__and3_1 c89 (.A(net65),
    .B(net64),
    .C(net1169),
    .X(net67));
 sky130_fd_sc_hd__and3_1 c90 (.A(net64),
    .B(net1169),
    .C(net913),
    .X(net68));
 sky130_fd_sc_hd__buf_1 c91 (.A(net867),
    .X(net69));
 sky130_fd_sc_hd__and3_1 c92 (.A(net63),
    .B(net68),
    .C(net1169),
    .X(net70));
 sky130_fd_sc_hd__and3_1 c93 (.A(net69),
    .B(net70),
    .C(net1169),
    .X(net71));
 sky130_fd_sc_hd__and3_1 c94 (.A(net68),
    .B(net65),
    .C(net1169),
    .X(net72));
 sky130_fd_sc_hd__a2111o_1 c95 (.A1(net67),
    .A2(net70),
    .B1(net69),
    .C1(net68),
    .D1(net1169),
    .X(net73));
 sky130_fd_sc_hd__mux4_1 c96 (.A0(net71),
    .A1(net64),
    .A2(net69),
    .A3(net73),
    .S0(net70),
    .S1(net1169),
    .X(net74));
 sky130_fd_sc_hd__mux4_1 c97 (.A0(net66),
    .A1(net69),
    .A2(net73),
    .A3(net1169),
    .S0(net68),
    .S1(net917),
    .X(net75));
 sky130_fd_sc_hd__sdfbbn_1 c98 (.CLK_N(clknet_leaf_44_clk),
    .D(net73),
    .RESET_B(net1171),
    .SCD(net71),
    .SCE(net72),
    .SET_B(net917),
    .Q(net77),
    .Q_N(net76));
 sky130_fd_sc_hd__mux4_1 c99 (.A0(net70),
    .A1(net73),
    .A2(net69),
    .A3(net1169),
    .S0(net913),
    .S1(net917),
    .X(net78));
 sky130_fd_sc_hd__a2111o_1 merge740 (.A1(net1163),
    .A2(net463),
    .B1(clknet_1_0__leaf_net465),
    .C1(net1177),
    .D1(net1035),
    .X(net761));
 sky130_fd_sc_hd__or4bb_1 merge741 (.A(net18),
    .B(net1166),
    .C_N(net1174),
    .D_N(net1235),
    .X(net762));
 sky130_fd_sc_hd__clkbuf_1 merge742 (.A(net793),
    .X(net763));
 sky130_fd_sc_hd__sdfbbn_1 merge743 (.CLK_N(clknet_leaf_42_clk),
    .D(clknet_1_1__leaf_net318),
    .RESET_B(net305),
    .SCE(net314),
    .SET_B(net995),
    .Q(net319),
    .Q_N(net764));
 sky130_fd_sc_hd__buf_1 merge744 (.A(net1125),
    .X(net766));
 sky130_fd_sc_hd__sdfrbp_1 merge745 (.CLK(clknet_leaf_46_clk),
    .D(net60),
    .RESET_B(net1170),
    .SCD(net86),
    .Q(net768),
    .Q_N(net767));
 sky130_fd_sc_hd__sdfrbp_2 merge746 (.CLK(clknet_leaf_21_clk),
    .D(net1267),
    .RESET_B(net712),
    .SCD(clknet_1_0__leaf_net1153),
    .Q(net713),
    .Q_N(net769));
 sky130_fd_sc_hd__clkbuf_1 merge747 (.A(net866),
    .X(net771));
 sky130_fd_sc_hd__clkbuf_1 merge748 (.A(net1120),
    .X(net772));
 sky130_fd_sc_hd__sdfrtn_1 merge749 (.CLK_N(clknet_leaf_10_clk),
    .D(clknet_1_0__leaf_net249),
    .RESET_B(clknet_1_0__leaf_net248),
    .SCD(net250),
    .SCE(clknet_1_0__leaf_net252),
    .Q(net773));
 sky130_fd_sc_hd__sdfrtp_1 merge750 (.CLK(clknet_leaf_10_clk),
    .D(net109),
    .RESET_B(net108),
    .SCD(net1208),
    .SCE(net826),
    .Q(net774));
 sky130_fd_sc_hd__clkbuf_1 merge751 (.A(net1125),
    .X(net775));
 sky130_fd_sc_hd__or4bb_1 merge752 (.A(clknet_1_1__leaf_net642),
    .B(clknet_1_1__leaf_net641),
    .C_N(net1182),
    .D_N(clknet_1_1__leaf_net548),
    .X(net776));
 sky130_fd_sc_hd__sdfrtp_1 merge753 (.CLK(clknet_leaf_25_clk),
    .D(clknet_1_1__leaf_net1154),
    .RESET_B(net741),
    .SCE(net1114),
    .Q(net739));
 sky130_fd_sc_hd__or4bb_1 merge754 (.A(net130),
    .B(net133),
    .C_N(net131),
    .D_N(net132),
    .X(net778));
 sky130_fd_sc_hd__sdfrtp_1 merge755 (.CLK(clknet_leaf_11_clk),
    .D(net393),
    .SCD(net395),
    .SCE(net930),
    .Q(net394));
 sky130_fd_sc_hd__sdfsbp_2 merge756 (.CLK(clknet_leaf_39_clk),
    .D(clknet_1_0__leaf_net105),
    .SCD(net214),
    .SET_B(clknet_1_1__leaf_net926),
    .Q(net224),
    .Q_N(net780));
 sky130_fd_sc_hd__or4bb_1 merge757 (.A(clknet_1_1__leaf_net618),
    .B(clknet_1_1__leaf_net619),
    .C_N(net1184),
    .D_N(net1090),
    .X(net782));
 sky130_fd_sc_hd__a2111o_1 merge758 (.A1(clknet_1_0__leaf_net596),
    .A2(clknet_1_0__leaf_net595),
    .B1(net597),
    .C1(net598),
    .D1(net1042),
    .X(net783));
 sky130_fd_sc_hd__or4bb_1 merge759 (.A(net1194),
    .B(net314),
    .C_N(net1188),
    .D_N(net305),
    .X(net784));
 sky130_fd_sc_hd__sdfsbp_1 merge760 (.CLK(clknet_leaf_8_clk),
    .D(net1210),
    .SCD(net393),
    .SCE(clknet_1_1__leaf_net157),
    .SET_B(clknet_1_1__leaf_net156),
    .Q(net786),
    .Q_N(net785));
 sky130_fd_sc_hd__or4bb_1 merge761 (.A(net1170),
    .B(net60),
    .C_N(net46),
    .D_N(net59),
    .X(net787));
 sky130_fd_sc_hd__mux4_1 merge762 (.A0(clknet_1_1__leaf_net1150),
    .A1(clknet_1_1__leaf_net507),
    .A2(net725),
    .A3(net714),
    .S0(net715),
    .S1(net1240),
    .X(net788));
 sky130_fd_sc_hd__mux4_1 merge763 (.A0(net322),
    .A1(net314),
    .A2(net1176),
    .A3(net320),
    .S0(clknet_1_1__leaf_net318),
    .S1(net1200),
    .X(net789));
 sky130_fd_sc_hd__sdfstp_1 merge764 (.CLK(clknet_leaf_14_clk),
    .D(clknet_1_0__leaf_net550),
    .SCD(clknet_1_0__leaf_net548),
    .SCE(clknet_1_1__leaf_net418),
    .SET_B(net419),
    .Q(net790));
 sky130_fd_sc_hd__sdfstp_2 merge765 (.CLK(clknet_leaf_27_clk),
    .D(net714),
    .SCD(net712),
    .SET_B(net1221),
    .Q(net715));
 sky130_fd_sc_hd__mux4_1 merge766 (.A0(net201),
    .A1(clknet_1_1__leaf_net205),
    .A2(clknet_1_1__leaf_net203),
    .A3(clknet_1_0__leaf_net1160),
    .S0(net511),
    .S1(clknet_1_0__leaf_net1150),
    .X(net792));
 sky130_fd_sc_hd__sdfstp_1 merge767 (.CLK(clknet_leaf_8_clk),
    .D(net1178),
    .SCD(net1165),
    .SCE(net269),
    .SET_B(net270),
    .Q(net793));
 sky130_fd_sc_hd__dfbbn_1 merge768 (.CLK_N(clknet_leaf_14_clk),
    .D(net527),
    .SET_B(net529),
    .Q(net795),
    .Q_N(net530));
 sky130_fd_sc_hd__sedfxbp_1 merge769 (.CLK(clknet_leaf_2_clk),
    .D(net109),
    .DE(net765),
    .SCD(net1207),
    .SCE(net113),
    .Q(net797),
    .Q_N(net796));
 sky130_fd_sc_hd__mux4_1 merge770 (.A0(net509),
    .A1(clknet_1_0__leaf_net1150),
    .A2(net370),
    .A3(net368),
    .S0(net1000),
    .S1(net1020),
    .X(net798));
 sky130_fd_sc_hd__mux4_1 merge771 (.A0(clknet_1_0__leaf_net689),
    .A1(net690),
    .A2(net1192),
    .A3(net527),
    .S0(net528),
    .S1(net1082),
    .X(net799));
 sky130_fd_sc_hd__mux4_1 merge772 (.A0(net41),
    .A1(net43),
    .A2(net1180),
    .A3(net23),
    .S0(net1166),
    .S1(net1174),
    .X(net800));
 sky130_fd_sc_hd__mux4_1 merge773 (.A0(net21),
    .A1(net22),
    .A2(net20),
    .A3(net275),
    .S0(net1178),
    .S1(net1165),
    .X(net801));
 sky130_fd_sc_hd__mux4_1 merge774 (.A0(net530),
    .A1(net532),
    .A2(net527),
    .A3(net274),
    .S0(net273),
    .S1(net271),
    .X(net802));
 sky130_fd_sc_hd__sdfbbp_1 merge775 (.CLK(clknet_leaf_17_clk),
    .D(net695),
    .RESET_B(clknet_1_0__leaf_net694),
    .SCD(net1172),
    .SCE(net582),
    .SET_B(net580),
    .Q(net804),
    .Q_N(net803));
 sky130_fd_sc_hd__sdfbbn_1 merge776 (.CLK_N(clknet_leaf_17_clk),
    .D(clknet_1_0__leaf_net694),
    .RESET_B(net695),
    .SCE(clknet_1_0__leaf_net574),
    .SET_B(net1238),
    .Q(net806),
    .Q_N(net805));
 sky130_fd_sc_hd__or4bb_1 merge777 (.A(net696),
    .B(net697),
    .C_N(clknet_1_1__leaf_net694),
    .D_N(net698),
    .X(net807));
 sky130_fd_sc_hd__mux4_1 merge778 (.A0(net153),
    .A1(net1165),
    .A2(net64),
    .A3(net60),
    .S0(net62),
    .S1(net1202),
    .X(net808));
 sky130_fd_sc_hd__dfrbp_1 merge779 (.CLK(clknet_leaf_40_clk),
    .D(net231),
    .RESET_B(net232),
    .Q(net810),
    .Q_N(net809));
 sky130_fd_sc_hd__dfrbp_1 merge780 (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1224),
    .Q(net812),
    .Q_N(net367));
 sky130_fd_sc_hd__dfrtn_1 merge781 (.CLK_N(clknet_leaf_5_clk),
    .D(net162),
    .RESET_B(net177),
    .Q(net813));
 sky130_fd_sc_hd__and2_0 merge782 (.A(net716),
    .B(net727),
    .X(net814));
 sky130_fd_sc_hd__dfrtp_1 merge783 (.CLK(clknet_leaf_36_clk),
    .D(net389),
    .RESET_B(net375),
    .Q(net815));
 sky130_fd_sc_hd__and2_0 merge784 (.A(net588),
    .B(net592),
    .X(net816));
 sky130_fd_sc_hd__dfrtp_1 merge785 (.CLK(clknet_leaf_13_clk),
    .D(net536),
    .RESET_B(net542),
    .Q(net817));
 sky130_fd_sc_hd__dfrtp_1 merge786 (.CLK(clknet_leaf_17_clk),
    .D(net573),
    .RESET_B(net561),
    .Q(net818));
 sky130_fd_sc_hd__dfsbp_1 merge787 (.CLK(clknet_leaf_17_clk),
    .D(net704),
    .SET_B(net708),
    .Q(net820),
    .Q_N(net819));
 sky130_fd_sc_hd__dfsbp_1 merge788 (.CLK(clknet_leaf_36_clk),
    .D(net515),
    .SET_B(net519),
    .Q(net822),
    .Q_N(net821));
 sky130_fd_sc_hd__dfstp_1 merge789 (.CLK(clknet_leaf_5_clk),
    .D(net300),
    .SET_B(net304),
    .Q(net823));
 sky130_fd_sc_hd__and2_0 merge790 (.A(net75),
    .B(net81),
    .X(net824));
 sky130_fd_sc_hd__dfstp_1 merge791 (.CLK(clknet_leaf_15_clk),
    .D(net432),
    .SET_B(net434),
    .Q(net825));
 sky130_fd_sc_hd__dfstp_1 merge792 (.CLK(clknet_leaf_10_clk),
    .D(net125),
    .SET_B(net112),
    .Q(net826));
 sky130_fd_sc_hd__dlrbn_1 merge793 (.D(net630),
    .GATE_N(clknet_leaf_32_clk),
    .RESET_B(net622),
    .Q(net828),
    .Q_N(net827));
 sky130_fd_sc_hd__and2_0 merge794 (.A(net8),
    .B(net15),
    .X(net829));
 sky130_fd_sc_hd__dlrbn_1 merge795 (.D(net460),
    .GATE_N(clknet_leaf_29_clk),
    .RESET_B(net784),
    .Q(net831),
    .Q_N(net830));
 sky130_fd_sc_hd__dlrbp_1 merge796 (.D(net152),
    .GATE(clknet_leaf_9_clk),
    .RESET_B(net778),
    .Q(net833),
    .Q_N(net832));
 sky130_fd_sc_hd__dlrbp_1 merge797 (.D(net494),
    .GATE(clknet_leaf_30_clk),
    .Q(net497),
    .Q_N(net834));
 sky130_fd_sc_hd__dlrtn_1 merge798 (.D(net259),
    .GATE_N(clknet_leaf_11_clk),
    .RESET_B(net265),
    .Q(net836));
 sky130_fd_sc_hd__dlrtn_1 merge799 (.D(net26),
    .GATE_N(clknet_leaf_1_clk),
    .Q(net29));
 sky130_fd_sc_hd__and2_0 merge800 (.A(net481),
    .B(net486),
    .X(net838));
 sky130_fd_sc_hd__dlrtn_1 merge801 (.D(net288),
    .GATE_N(clknet_leaf_7_clk),
    .Q(net292));
 sky130_fd_sc_hd__dlrtp_1 merge802 (.D(net405),
    .GATE(clknet_leaf_12_clk),
    .RESET_B(net406),
    .Q(net840));
 sky130_fd_sc_hd__dlrtp_1 merge803 (.D(net99),
    .GATE(clknet_leaf_45_clk),
    .RESET_B(net104),
    .Q(net841));
 sky130_fd_sc_hd__dlrtp_1 merge804 (.D(net61),
    .GATE(clknet_leaf_47_clk),
    .RESET_B(net49),
    .Q(net842));
 sky130_fd_sc_hd__edfxbp_1 merge805 (.CLK(clknet_leaf_4_clk),
    .DE(net187),
    .Q(net844),
    .Q_N(net189));
 sky130_fd_sc_hd__edfxtp_1 merge806 (.CLK(clknet_leaf_23_clk),
    .D(net753),
    .Q(net845));
 sky130_fd_sc_hd__sdlclkp_1 merge807 (.CLK(clknet_leaf_41_clk),
    .GATE(net209),
    .SCE(net217),
    .GCLK(net846));
 sky130_fd_sc_hd__and2_0 merge808 (.A(net654),
    .B(net660),
    .X(net847));
 sky130_fd_sc_hd__sdlclkp_2 merge809 (.CLK(clknet_leaf_31_clk),
    .GATE(net617),
    .SCE(net607),
    .GCLK(net848));
 sky130_fd_sc_hd__and2_0 merge810 (.A(net324),
    .B(net336),
    .X(net849));
 sky130_fd_sc_hd__and2_0 merge811 (.A(net679),
    .B(net682),
    .X(net850));
 sky130_fd_sc_hd__and2_0 merge812 (.A(net315),
    .B(net83),
    .X(net851));
 sky130_fd_sc_hd__and2_0 merge813 (.A(net16),
    .B(net178),
    .X(net852));
 sky130_fd_sc_hd__and2_0 merge814 (.A(net82),
    .B(net235),
    .X(net853));
 sky130_fd_sc_hd__and2_0 merge815 (.A(net526),
    .B(net245),
    .X(net854));
 sky130_fd_sc_hd__sdlclkp_4 merge816 (.CLK(clknet_leaf_2_clk),
    .GATE(net829),
    .SCE(net119),
    .GCLK(net855));
 sky130_fd_sc_hd__dfrbp_1 merge817 (.CLK(clknet_leaf_7_clk),
    .D(net439),
    .RESET_B(net268),
    .Q(net857),
    .Q_N(net856));
 sky130_fd_sc_hd__dfrbp_1 merge818 (.CLK(clknet_leaf_27_clk),
    .D(net594),
    .RESET_B(net728),
    .Q(net859),
    .Q_N(net858));
 sky130_fd_sc_hd__and2_0 merge819 (.A(net759),
    .B(net734),
    .X(net860));
 sky130_fd_sc_hd__dfrtn_1 merge820 (.CLK_N(clknet_leaf_36_clk),
    .D(net520),
    .RESET_B(net388),
    .Q(net861));
 sky130_fd_sc_hd__and2_0 merge821 (.A(net313),
    .B(net317),
    .X(net862));
 sky130_fd_sc_hd__and2_0 merge822 (.A(net688),
    .B(net666),
    .X(net863));
 sky130_fd_sc_hd__dfrtp_1 merge823 (.CLK(clknet_leaf_25_clk),
    .D(net757),
    .RESET_B(net632),
    .Q(net864));
 sky130_fd_sc_hd__dfrtp_1 merge824 (.CLK(clknet_leaf_3_clk),
    .D(net39),
    .RESET_B(net762),
    .Q(net865));
 sky130_fd_sc_hd__dfrtp_1 merge825 (.CLK(clknet_leaf_39_clk),
    .D(net244),
    .RESET_B(net787),
    .Q(net866));
 sky130_fd_sc_hd__dfsbp_1 merge826 (.CLK(clknet_leaf_8_clk),
    .D(net267),
    .SET_B(net808),
    .Q(net868),
    .Q_N(net867));
 sky130_fd_sc_hd__dfsbp_1 merge827 (.CLK(clknet_leaf_23_clk),
    .D(net733),
    .SET_B(net687),
    .Q(net870),
    .Q_N(net869));
 sky130_fd_sc_hd__dfstp_1 merge828 (.CLK(clknet_leaf_16_clk),
    .SET_B(net437),
    .Q(net438));
 sky130_fd_sc_hd__dfstp_1 merge829 (.CLK(clknet_leaf_21_clk),
    .D(net776),
    .SET_B(net850),
    .Q(net872));
 sky130_fd_sc_hd__dfstp_2 merge830 (.CLK(clknet_leaf_16_clk),
    .D(net277),
    .SET_B(net862),
    .Q(net873));
 sky130_fd_sc_hd__dlrbn_1 merge831 (.D(net782),
    .GATE_N(clknet_leaf_26_clk),
    .RESET_B(net638),
    .Q(net875),
    .Q_N(net874));
 sky130_fd_sc_hd__dlrbn_1 merge832 (.D(net847),
    .GATE_N(clknet_leaf_17_clk),
    .RESET_B(net807),
    .Q(net877),
    .Q_N(net876));
 sky130_fd_sc_hd__dlrbp_1 merge833 (.D(net838),
    .GATE(clknet_leaf_30_clk),
    .RESET_B(net508),
    .Q(net879),
    .Q_N(net878));
 sky130_fd_sc_hd__dlrbp_1 merge834 (.D(net849),
    .GATE(clknet_leaf_43_clk),
    .RESET_B(net852),
    .Q(net881),
    .Q_N(net880));
 sky130_fd_sc_hd__dlrtn_1 merge835 (.D(net863),
    .GATE_N(clknet_leaf_20_clk),
    .RESET_B(net677),
    .Q(net882));
 sky130_fd_sc_hd__dlrtn_1 merge836 (.D(net625),
    .GATE_N(clknet_leaf_26_clk),
    .RESET_B(net816),
    .Q(net883));
 sky130_fd_sc_hd__dlrtn_1 merge837 (.D(net824),
    .GATE_N(clknet_leaf_40_clk),
    .RESET_B(net853),
    .Q(net884));
 sky130_fd_sc_hd__dlrtp_1 merge838 (.D(net484),
    .GATE(clknet_leaf_30_clk),
    .RESET_B(net854),
    .Q(net1149));
 sky130_fd_sc_hd__dlrtp_1 merge839 (.D(net572),
    .GATE(clknet_leaf_17_clk),
    .RESET_B(net783),
    .Q(net885));
 sky130_fd_sc_hd__dlrtp_1 merge840 (.D(net628),
    .GATE(clknet_leaf_33_clk),
    .Q(net886));
 sky130_fd_sc_hd__edfxbp_1 merge841 (.CLK(clknet_leaf_21_clk),
    .D(net675),
    .DE(net814),
    .Q(net888),
    .Q_N(net887));
 sky130_fd_sc_hd__edfxtp_1 merge842 (.CLK(clknet_leaf_0_clk),
    .D(net53),
    .DE(net30),
    .Q(net889));
 sky130_fd_sc_hd__sdlclkp_1 merge843 (.CLK(clknet_leaf_5_clk),
    .GATE(net176),
    .SCE(net761),
    .GCLK(net890));
 sky130_fd_sc_hd__sdlclkp_2 merge844 (.CLK(clknet_leaf_29_clk),
    .GATE(net851),
    .SCE(net593),
    .GCLK(net891));
 sky130_fd_sc_hd__sdlclkp_4 merge845 (.CLK(clknet_leaf_31_clk),
    .GATE(net610),
    .SCE(net506),
    .GCLK(net892));
 sky130_fd_sc_hd__dfrbp_1 merge846 (.CLK(clknet_leaf_35_clk),
    .D(net792),
    .RESET_B(net387),
    .Q(net894),
    .Q_N(net893));
 sky130_fd_sc_hd__dfrbp_1 merge847 (.CLK(clknet_leaf_27_clk),
    .D(net709),
    .RESET_B(net860),
    .Q(net896),
    .Q_N(net895));
 sky130_fd_sc_hd__dlxbn_1 s1000 (.D(net635),
    .GATE_N(clknet_leaf_26_clk),
    .Q(net1155),
    .Q_N(net1094));
 sky130_fd_sc_hd__dlxbn_1 s1001 (.D(net637),
    .GATE_N(clknet_leaf_25_clk),
    .Q(net1096),
    .Q_N(net1095));
 sky130_fd_sc_hd__dlxbp_1 s1002 (.D(net640),
    .GATE(clknet_leaf_33_clk),
    .Q(net1151),
    .Q_N(net1152));
 sky130_fd_sc_hd__dlxtn_1 s1003 (.D(net649),
    .GATE_N(clknet_leaf_18_clk),
    .Q(net1097));
 sky130_fd_sc_hd__dlxtn_1 s1004 (.D(net657),
    .GATE_N(clknet_leaf_19_clk),
    .Q(net1098));
 sky130_fd_sc_hd__dlxtn_1 s1005 (.D(net658),
    .GATE_N(clknet_leaf_19_clk),
    .Q(net1099));
 sky130_fd_sc_hd__dlxtp_1 s1006 (.D(net659),
    .GATE(clknet_leaf_19_clk),
    .Q(net1100));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s1007 (.D(net661),
    .SLEEP_B(clknet_leaf_20_clk),
    .Q(net1101));
 sky130_fd_sc_hd__dfxbp_1 s1008 (.CLK(clknet_leaf_20_clk),
    .D(net674),
    .Q(net1103),
    .Q_N(net1102));
 sky130_fd_sc_hd__dfxbp_1 s1009 (.CLK(clknet_leaf_20_clk),
    .D(net676),
    .Q(net1105),
    .Q_N(net1104));
 sky130_fd_sc_hd__dfxtp_1 s1010 (.CLK(clknet_leaf_22_clk),
    .D(net678),
    .Q(net1106));
 sky130_fd_sc_hd__dfxtp_2 s1011 (.CLK(clknet_leaf_22_clk),
    .D(net680),
    .Q(net1107));
 sky130_fd_sc_hd__dfxtp_1 s1012 (.CLK(clknet_leaf_22_clk),
    .D(net683),
    .Q(net1108));
 sky130_fd_sc_hd__dlclkp_1 s1013 (.CLK(clknet_leaf_21_clk),
    .GATE(net684),
    .GCLK(net1109));
 sky130_fd_sc_hd__dlclkp_2 s1014 (.CLK(clknet_leaf_21_clk),
    .GATE(net685),
    .GCLK(net1110));
 sky130_fd_sc_hd__dlclkp_4 s1015 (.CLK(clknet_leaf_22_clk),
    .GATE(net686),
    .GCLK(net1111));
 sky130_fd_sc_hd__dlxbn_1 s1016 (.D(net732),
    .GATE_N(clknet_leaf_23_clk),
    .Q(net1113),
    .Q_N(net1112));
 sky130_fd_sc_hd__dlxbn_1 s1017 (.D(net735),
    .GATE_N(clknet_leaf_23_clk),
    .Q(net1115),
    .Q_N(net1114));
 sky130_fd_sc_hd__dlxbp_1 s1018 (.D(net750),
    .GATE(clknet_leaf_23_clk),
    .Q(net1117),
    .Q_N(net1116));
 sky130_fd_sc_hd__dlxtn_1 s1019 (.D(net752),
    .GATE_N(clknet_leaf_23_clk),
    .Q(net1118));
 sky130_fd_sc_hd__dlxtn_1 s1020 (.D(net755),
    .GATE_N(clknet_leaf_23_clk),
    .Q(net1119));
 sky130_fd_sc_hd__dlxtn_1 s1021 (.D(net756),
    .GATE_N(clknet_leaf_24_clk),
    .Q(net1159));
 sky130_fd_sc_hd__dlxtp_1 s1022 (.D(net760),
    .GATE(clknet_leaf_25_clk),
    .Q(net1158));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s1023 (.D(net788),
    .SLEEP_B(clknet_leaf_32_clk),
    .Q(net1120));
 sky130_fd_sc_hd__dfxbp_1 s1024 (.CLK(clknet_leaf_42_clk),
    .D(net789),
    .Q(net1122),
    .Q_N(net1121));
 sky130_fd_sc_hd__dfxbp_1 s1025 (.CLK(clknet_leaf_35_clk),
    .D(net798),
    .Q(net1124),
    .Q_N(net1123));
 sky130_fd_sc_hd__dfxtp_1 s1026 (.CLK(clknet_leaf_17_clk),
    .D(net799),
    .Q(net1125));
 sky130_fd_sc_hd__dfxtp_1 s1027 (.CLK(clknet_leaf_0_clk),
    .D(net800),
    .Q(net1126));
 sky130_fd_sc_hd__dfxtp_1 s1028 (.CLK(clknet_leaf_3_clk),
    .D(net801),
    .Q(net1127));
 sky130_fd_sc_hd__dlclkp_1 s1029 (.CLK(clknet_leaf_15_clk),
    .GATE(net802),
    .GCLK(net1128));
 sky130_fd_sc_hd__dfxbp_1 s848 (.CLK(clknet_leaf_1_clk),
    .D(net6),
    .Q(net898),
    .Q_N(net897));
 sky130_fd_sc_hd__dfxbp_1 s849 (.CLK(clknet_leaf_1_clk),
    .D(net7),
    .Q(net900),
    .Q_N(net899));
 sky130_fd_sc_hd__dfxtp_1 s850 (.CLK(clknet_leaf_1_clk),
    .D(net10),
    .Q(net901));
 sky130_fd_sc_hd__dfxtp_1 s851 (.CLK(clknet_leaf_1_clk),
    .D(net13),
    .Q(net902));
 sky130_fd_sc_hd__dfxtp_1 s852 (.CLK(clknet_leaf_2_clk),
    .D(net17),
    .Q(net903));
 sky130_fd_sc_hd__dlclkp_1 s853 (.CLK(clknet_leaf_0_clk),
    .GATE(net31),
    .GCLK(net904));
 sky130_fd_sc_hd__dlclkp_2 s854 (.CLK(clknet_leaf_3_clk),
    .GATE(net32),
    .GCLK(net905));
 sky130_fd_sc_hd__dlclkp_4 s855 (.CLK(clknet_leaf_0_clk),
    .GATE(net33),
    .GCLK(net906));
 sky130_fd_sc_hd__dlxbn_2 s856 (.D(net34),
    .GATE_N(clknet_leaf_0_clk),
    .Q(net908),
    .Q_N(net907));
 sky130_fd_sc_hd__dlxbn_1 s857 (.D(net36),
    .GATE_N(clknet_leaf_3_clk),
    .Q(net910),
    .Q_N(net909));
 sky130_fd_sc_hd__dlxbp_1 s858 (.D(net51),
    .GATE(clknet_leaf_48_clk),
    .Q(net912),
    .Q_N(net911));
 sky130_fd_sc_hd__dlxtn_2 s859 (.D(net52),
    .GATE_N(clknet_leaf_47_clk),
    .Q(net913));
 sky130_fd_sc_hd__dlxtn_1 s860 (.D(net55),
    .GATE_N(clknet_leaf_48_clk),
    .Q(net914));
 sky130_fd_sc_hd__dlxtn_1 s861 (.D(net56),
    .GATE_N(clknet_leaf_48_clk),
    .Q(net915));
 sky130_fd_sc_hd__dlxtp_1 s862 (.D(net57),
    .GATE(clknet_leaf_48_clk),
    .Q(net916));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s863 (.D(net74),
    .SLEEP_B(clknet_leaf_46_clk),
    .Q(net917));
 sky130_fd_sc_hd__dfxbp_1 s864 (.CLK(clknet_leaf_44_clk),
    .D(net78),
    .Q(net919),
    .Q_N(net918));
 sky130_fd_sc_hd__dfxbp_1 s865 (.CLK(clknet_leaf_45_clk),
    .D(net79),
    .Q(net921),
    .Q_N(net920));
 sky130_fd_sc_hd__dfxtp_1 s866 (.CLK(clknet_leaf_46_clk),
    .D(net92),
    .Q(net922));
 sky130_fd_sc_hd__dfxtp_1 s867 (.CLK(clknet_leaf_45_clk),
    .D(net101),
    .Q(net923));
 sky130_fd_sc_hd__dfxtp_1 s868 (.CLK(clknet_leaf_45_clk),
    .D(net102),
    .Q(net924));
 sky130_fd_sc_hd__dlclkp_1 s869 (.CLK(clknet_leaf_39_clk),
    .GATE(net103),
    .GCLK(net925));
 sky130_fd_sc_hd__dlclkp_2 s870 (.CLK(clknet_leaf_39_clk),
    .GATE(net106),
    .GCLK(net926));
 sky130_fd_sc_hd__dlclkp_4 s871 (.CLK(clknet_leaf_9_clk),
    .GATE(net124),
    .GCLK(net927));
 sky130_fd_sc_hd__dlxbn_1 s872 (.D(net126),
    .GATE_N(clknet_leaf_10_clk),
    .Q(net929),
    .Q_N(net928));
 sky130_fd_sc_hd__dlxbn_1 s873 (.D(net128),
    .GATE_N(clknet_leaf_10_clk),
    .Q(net931),
    .Q_N(net930));
 sky130_fd_sc_hd__dlxbp_1 s874 (.D(net129),
    .GATE(clknet_leaf_10_clk),
    .Q(net933),
    .Q_N(net932));
 sky130_fd_sc_hd__dlxtn_1 s875 (.D(net144),
    .GATE_N(clknet_leaf_2_clk),
    .Q(net934));
 sky130_fd_sc_hd__dlxtn_1 s876 (.D(net145),
    .GATE_N(clknet_leaf_2_clk),
    .Q(net935));
 sky130_fd_sc_hd__dlxtn_1 s877 (.D(net146),
    .GATE_N(clknet_leaf_8_clk),
    .Q(net936));
 sky130_fd_sc_hd__dlxtp_1 s878 (.D(net149),
    .GATE(clknet_leaf_9_clk),
    .Q(net937));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s879 (.D(net150),
    .SLEEP_B(clknet_leaf_9_clk),
    .Q(net938));
 sky130_fd_sc_hd__dfxbp_1 s880 (.CLK(clknet_leaf_9_clk),
    .D(net151),
    .Q(net940),
    .Q_N(net939));
 sky130_fd_sc_hd__dfxbp_1 s881 (.CLK(clknet_leaf_4_clk),
    .D(net167),
    .Q(net942),
    .Q_N(net941));
 sky130_fd_sc_hd__dfxtp_1 s882 (.CLK(clknet_leaf_4_clk),
    .D(net168),
    .Q(net943));
 sky130_fd_sc_hd__dfxtp_1 s883 (.CLK(clknet_leaf_4_clk),
    .D(net169),
    .Q(net944));
 sky130_fd_sc_hd__dfxtp_1 s884 (.CLK(clknet_leaf_5_clk),
    .D(net170),
    .Q(net945));
 sky130_fd_sc_hd__dlclkp_1 s885 (.CLK(clknet_leaf_5_clk),
    .GATE(net172),
    .GCLK(net946));
 sky130_fd_sc_hd__dlclkp_2 s886 (.CLK(clknet_leaf_43_clk),
    .GATE(net173),
    .GCLK(net947));
 sky130_fd_sc_hd__dlclkp_4 s887 (.CLK(clknet_leaf_43_clk),
    .GATE(net174),
    .GCLK(net948));
 sky130_fd_sc_hd__dlxbn_1 s888 (.D(net175),
    .GATE_N(clknet_leaf_5_clk),
    .Q(net950),
    .Q_N(net949));
 sky130_fd_sc_hd__dlxbn_1 s889 (.D(net186),
    .GATE_N(clknet_leaf_47_clk),
    .Q(net952),
    .Q_N(net951));
 sky130_fd_sc_hd__dlxbp_1 s890 (.D(net188),
    .GATE(clknet_leaf_44_clk),
    .Q(net954),
    .Q_N(net953));
 sky130_fd_sc_hd__dlxtn_1 s891 (.D(net190),
    .GATE_N(clknet_leaf_44_clk),
    .Q(net955));
 sky130_fd_sc_hd__dlxtn_1 s892 (.D(net191),
    .GATE_N(clknet_leaf_44_clk),
    .Q(net956));
 sky130_fd_sc_hd__dlxtn_1 s893 (.D(net192),
    .GATE_N(clknet_leaf_44_clk),
    .Q(net957));
 sky130_fd_sc_hd__dlxtp_1 s894 (.D(net193),
    .GATE(clknet_leaf_44_clk),
    .Q(net958));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s895 (.D(net194),
    .SLEEP_B(clknet_leaf_43_clk),
    .Q(net959));
 sky130_fd_sc_hd__dfxbp_1 s896 (.CLK(clknet_leaf_44_clk),
    .D(net196),
    .Q(net961),
    .Q_N(net960));
 sky130_fd_sc_hd__dfxbp_1 s897 (.CLK(clknet_leaf_43_clk),
    .D(net197),
    .Q(net963),
    .Q_N(net962));
 sky130_fd_sc_hd__dfxtp_1 s898 (.CLK(clknet_leaf_43_clk),
    .D(net198),
    .Q(net964));
 sky130_fd_sc_hd__dfxtp_1 s899 (.CLK(clknet_leaf_40_clk),
    .D(net218),
    .Q(net965));
 sky130_fd_sc_hd__dfxtp_1 s900 (.CLK(clknet_leaf_40_clk),
    .D(net219),
    .Q(net966));
 sky130_fd_sc_hd__dlclkp_1 s901 (.CLK(clknet_leaf_40_clk),
    .GATE(net221),
    .GCLK(net967));
 sky130_fd_sc_hd__dlclkp_2 s902 (.CLK(clknet_leaf_40_clk),
    .GATE(net222),
    .GCLK(net968));
 sky130_fd_sc_hd__dlclkp_4 s903 (.CLK(clknet_leaf_40_clk),
    .GATE(net223),
    .GCLK(net969));
 sky130_fd_sc_hd__dlxbn_1 s904 (.D(net236),
    .GATE_N(clknet_leaf_39_clk),
    .Q(net971),
    .Q_N(net970));
 sky130_fd_sc_hd__dlxbn_1 s905 (.D(net237),
    .GATE_N(clknet_leaf_39_clk),
    .Q(net973),
    .Q_N(net972));
 sky130_fd_sc_hd__dlxbp_1 s906 (.D(net239),
    .GATE(clknet_leaf_38_clk),
    .Q(net975),
    .Q_N(net974));
 sky130_fd_sc_hd__dlxtn_1 s907 (.D(net240),
    .GATE_N(clknet_leaf_39_clk),
    .Q(net976));
 sky130_fd_sc_hd__dlxtn_1 s908 (.D(net241),
    .GATE_N(clknet_leaf_38_clk),
    .Q(net977));
 sky130_fd_sc_hd__dlxtn_1 s909 (.D(net246),
    .GATE_N(clknet_leaf_35_clk),
    .Q(net978));
 sky130_fd_sc_hd__dlxtp_1 s910 (.D(net258),
    .GATE(clknet_leaf_11_clk),
    .Q(net979));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s911 (.D(net261),
    .SLEEP_B(clknet_leaf_11_clk),
    .Q(net980));
 sky130_fd_sc_hd__dfxbp_1 s912 (.CLK(clknet_leaf_11_clk),
    .D(net262),
    .Q(net982),
    .Q_N(net981));
 sky130_fd_sc_hd__dfxbp_1 s913 (.CLK(clknet_leaf_11_clk),
    .D(net263),
    .Q(net984),
    .Q_N(net983));
 sky130_fd_sc_hd__dfxtp_1 s914 (.CLK(clknet_leaf_11_clk),
    .D(net264),
    .Q(net985));
 sky130_fd_sc_hd__dfxtp_1 s915 (.CLK(clknet_leaf_7_clk),
    .D(net282),
    .Q(net986));
 sky130_fd_sc_hd__dfxtp_1 s916 (.CLK(clknet_leaf_7_clk),
    .D(net285),
    .Q(net987));
 sky130_fd_sc_hd__dlclkp_1 s917 (.CLK(clknet_leaf_7_clk),
    .GATE(net286),
    .GCLK(net988));
 sky130_fd_sc_hd__dlclkp_2 s918 (.CLK(clknet_leaf_7_clk),
    .GATE(net287),
    .GCLK(net989));
 sky130_fd_sc_hd__dlclkp_4 s919 (.CLK(clknet_leaf_15_clk),
    .GATE(net289),
    .GCLK(net990));
 sky130_fd_sc_hd__dlxbn_1 s920 (.D(net291),
    .GATE_N(clknet_leaf_7_clk),
    .Q(net992),
    .Q_N(net991));
 sky130_fd_sc_hd__dlxbn_1 s921 (.D(net301),
    .GATE_N(clknet_leaf_6_clk),
    .Q(net994),
    .Q_N(net993));
 sky130_fd_sc_hd__dlxbp_1 s922 (.D(net316),
    .GATE(clknet_leaf_6_clk),
    .Q(net996),
    .Q_N(net995));
 sky130_fd_sc_hd__dlxtn_1 s923 (.D(net335),
    .GATE_N(clknet_leaf_42_clk),
    .Q(net997));
 sky130_fd_sc_hd__dlxtn_1 s924 (.D(net338),
    .GATE_N(clknet_leaf_42_clk),
    .Q(net998));
 sky130_fd_sc_hd__dlxtn_1 s925 (.D(net340),
    .GATE_N(clknet_leaf_42_clk),
    .Q(net999));
 sky130_fd_sc_hd__dlxtp_1 s926 (.D(net354),
    .GATE(clknet_leaf_41_clk),
    .Q(net1000));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s927 (.D(net357),
    .SLEEP_B(clknet_leaf_41_clk),
    .Q(net1001));
 sky130_fd_sc_hd__dfxbp_1 s928 (.CLK(clknet_leaf_38_clk),
    .D(net361),
    .Q(net1003),
    .Q_N(net1002));
 sky130_fd_sc_hd__dfxbp_1 s929 (.CLK(clknet_leaf_38_clk),
    .D(net362),
    .Q(net1005),
    .Q_N(net1004));
 sky130_fd_sc_hd__dfxtp_1 s930 (.CLK(clknet_leaf_38_clk),
    .D(net364),
    .Q(net1006));
 sky130_fd_sc_hd__dfxtp_1 s931 (.CLK(clknet_leaf_38_clk),
    .D(net365),
    .Q(net1007));
 sky130_fd_sc_hd__dfxtp_2 s932 (.CLK(clknet_leaf_37_clk),
    .D(net376),
    .Q(net1008));
 sky130_fd_sc_hd__dlclkp_1 s933 (.CLK(clknet_leaf_37_clk),
    .GATE(net377),
    .GCLK(net1009));
 sky130_fd_sc_hd__dlclkp_2 s934 (.CLK(clknet_leaf_37_clk),
    .GATE(net378),
    .GCLK(net1010));
 sky130_fd_sc_hd__dlclkp_4 s935 (.CLK(clknet_leaf_37_clk),
    .GATE(net379),
    .GCLK(net1011));
 sky130_fd_sc_hd__dlxbn_1 s936 (.D(net380),
    .GATE_N(clknet_leaf_37_clk),
    .Q(net1013),
    .Q_N(net1012));
 sky130_fd_sc_hd__dlxbn_1 s937 (.D(net382),
    .GATE_N(clknet_leaf_37_clk),
    .Q(net1015),
    .Q_N(net1014));
 sky130_fd_sc_hd__dlxbp_1 s938 (.D(net383),
    .GATE(clknet_leaf_36_clk),
    .Q(net1017),
    .Q_N(net1016));
 sky130_fd_sc_hd__dlxtn_1 s939 (.D(net384),
    .GATE_N(clknet_leaf_37_clk),
    .Q(net1018));
 sky130_fd_sc_hd__dlxtn_1 s940 (.D(net386),
    .GATE_N(clknet_leaf_36_clk),
    .Q(net1019));
 sky130_fd_sc_hd__dlxtn_2 s941 (.D(net390),
    .GATE_N(clknet_leaf_36_clk),
    .Q(net1020));
 sky130_fd_sc_hd__dlxtp_1 s942 (.D(net409),
    .GATE(clknet_leaf_12_clk),
    .Q(net1021));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s943 (.D(net410),
    .SLEEP_B(clknet_leaf_12_clk),
    .Q(net1022));
 sky130_fd_sc_hd__dfxbp_1 s944 (.CLK(clknet_leaf_14_clk),
    .D(net411),
    .Q(net1024),
    .Q_N(net1023));
 sky130_fd_sc_hd__dfxbp_1 s945 (.CLK(clknet_leaf_14_clk),
    .D(net412),
    .Q(net1026),
    .Q_N(net1025));
 sky130_fd_sc_hd__dfxtp_1 s946 (.CLK(clknet_leaf_16_clk),
    .D(net429),
    .Q(net1027));
 sky130_fd_sc_hd__dfxtp_1 s947 (.CLK(clknet_leaf_16_clk),
    .D(net433),
    .Q(net1028));
 sky130_fd_sc_hd__dfxtp_1 s948 (.CLK(clknet_leaf_16_clk),
    .D(net451),
    .Q(net1029));
 sky130_fd_sc_hd__dlclkp_1 s949 (.CLK(clknet_leaf_16_clk),
    .GATE(net452),
    .GCLK(net1030));
 sky130_fd_sc_hd__dlclkp_2 s950 (.CLK(clknet_leaf_16_clk),
    .GATE(net453),
    .GCLK(net1031));
 sky130_fd_sc_hd__dlclkp_4 s951 (.CLK(clknet_leaf_29_clk),
    .GATE(net454),
    .GCLK(net1032));
 sky130_fd_sc_hd__dlxbn_1 s952 (.D(net456),
    .GATE_N(clknet_leaf_28_clk),
    .Q(net1034),
    .Q_N(net1033));
 sky130_fd_sc_hd__dlxbn_2 s953 (.D(net461),
    .GATE_N(clknet_leaf_29_clk),
    .Q(net1036),
    .Q_N(net1035));
 sky130_fd_sc_hd__dlxbp_1 s954 (.D(net470),
    .GATE(clknet_leaf_42_clk),
    .Q(net1038),
    .Q_N(net1037));
 sky130_fd_sc_hd__dlxtn_1 s955 (.D(net475),
    .GATE_N(clknet_leaf_41_clk),
    .Q(net1039));
 sky130_fd_sc_hd__dlxtn_1 s956 (.D(net478),
    .GATE_N(clknet_leaf_29_clk),
    .Q(net1040));
 sky130_fd_sc_hd__dlxtn_1 s957 (.D(net480),
    .GATE_N(clknet_leaf_30_clk),
    .Q(net1041));
 sky130_fd_sc_hd__dlxtp_1 s958 (.D(net485),
    .GATE(clknet_leaf_41_clk),
    .Q(net1042));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s959 (.D(net493),
    .SLEEP_B(clknet_leaf_30_clk),
    .Q(net1043));
 sky130_fd_sc_hd__dfxbp_1 s960 (.CLK(clknet_leaf_31_clk),
    .D(net495),
    .Q(net1045),
    .Q_N(net1044));
 sky130_fd_sc_hd__dfxbp_1 s961 (.CLK(clknet_leaf_35_clk),
    .D(net496),
    .Q(net1047),
    .Q_N(net1046));
 sky130_fd_sc_hd__dfxtp_2 s962 (.CLK(clknet_leaf_34_clk),
    .D(net498),
    .Q(net1048));
 sky130_fd_sc_hd__dfxtp_1 s963 (.CLK(clknet_leaf_34_clk),
    .D(net500),
    .Q(net1049));
 sky130_fd_sc_hd__dfxtp_1 s964 (.CLK(clknet_leaf_32_clk),
    .D(net501),
    .Q(net1156));
 sky130_fd_sc_hd__dlclkp_1 s965 (.CLK(clknet_leaf_34_clk),
    .GATE(net502),
    .GCLK(net1050));
 sky130_fd_sc_hd__dlclkp_2 s966 (.CLK(clknet_leaf_34_clk),
    .GATE(net504),
    .GCLK(net1051));
 sky130_fd_sc_hd__dlclkp_4 s967 (.CLK(clknet_leaf_31_clk),
    .GATE(net505),
    .GCLK(net1052));
 sky130_fd_sc_hd__dlxbn_1 s968 (.D(net514),
    .GATE_N(clknet_leaf_34_clk),
    .Q(net1054),
    .Q_N(net1053));
 sky130_fd_sc_hd__dlxbn_1 s969 (.D(net516),
    .GATE_N(clknet_leaf_34_clk),
    .Q(net1056),
    .Q_N(net1055));
 sky130_fd_sc_hd__dlxbp_1 s970 (.D(net521),
    .GATE(clknet_leaf_33_clk),
    .Q(net1058),
    .Q_N(net1057));
 sky130_fd_sc_hd__dlxtn_1 s971 (.D(net522),
    .GATE_N(clknet_leaf_33_clk),
    .Q(net1059));
 sky130_fd_sc_hd__dlxtn_1 s972 (.D(net525),
    .GATE_N(clknet_leaf_33_clk),
    .Q(net1148));
 sky130_fd_sc_hd__dlxtn_1 s973 (.D(net540),
    .GATE_N(clknet_leaf_13_clk),
    .Q(net1060));
 sky130_fd_sc_hd__dlxtp_1 s974 (.D(net541),
    .GATE(clknet_leaf_13_clk),
    .Q(net1061));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s975 (.D(net543),
    .SLEEP_B(clknet_leaf_13_clk),
    .Q(net1062));
 sky130_fd_sc_hd__dfxbp_1 s976 (.CLK(clknet_leaf_13_clk),
    .D(net544),
    .Q(net1064),
    .Q_N(net1063));
 sky130_fd_sc_hd__dfxbp_1 s977 (.CLK(clknet_leaf_13_clk),
    .D(net545),
    .Q(net1066),
    .Q_N(net1065));
 sky130_fd_sc_hd__dfxtp_1 s978 (.CLK(clknet_leaf_13_clk),
    .D(net546),
    .Q(net1067));
 sky130_fd_sc_hd__dfxtp_1 s979 (.CLK(clknet_leaf_13_clk),
    .D(net547),
    .Q(net1068));
 sky130_fd_sc_hd__dfxtp_1 s980 (.CLK(clknet_leaf_16_clk),
    .D(net564),
    .Q(net1069));
 sky130_fd_sc_hd__dlclkp_1 s981 (.CLK(clknet_leaf_18_clk),
    .GATE(net565),
    .GCLK(net1070));
 sky130_fd_sc_hd__dlclkp_2 s982 (.CLK(clknet_leaf_18_clk),
    .GATE(net568),
    .GCLK(net1071));
 sky130_fd_sc_hd__dlclkp_4 s983 (.CLK(clknet_leaf_17_clk),
    .GATE(net569),
    .GCLK(net1072));
 sky130_fd_sc_hd__dlxbn_1 s984 (.D(net571),
    .GATE_N(clknet_leaf_17_clk),
    .Q(net1074),
    .Q_N(net1073));
 sky130_fd_sc_hd__dlxbn_1 s985 (.D(net584),
    .GATE_N(clknet_leaf_27_clk),
    .Q(net1076),
    .Q_N(net1075));
 sky130_fd_sc_hd__dlxbp_1 s986 (.D(net586),
    .GATE(clknet_leaf_28_clk),
    .Q(net1078),
    .Q_N(net1077));
 sky130_fd_sc_hd__dlxtn_1 s987 (.D(net587),
    .GATE_N(clknet_leaf_28_clk),
    .Q(net1079));
 sky130_fd_sc_hd__dlxtn_4 s988 (.D(net589),
    .GATE_N(clknet_leaf_27_clk),
    .Q(net1080));
 sky130_fd_sc_hd__dlxtn_1 s989 (.D(net590),
    .GATE_N(clknet_leaf_27_clk),
    .Q(net1081));
 sky130_fd_sc_hd__dlxtp_1 s990 (.D(net591),
    .GATE(clknet_leaf_27_clk),
    .Q(net1082));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s991 (.D(net603),
    .SLEEP_B(clknet_leaf_28_clk),
    .Q(net1083));
 sky130_fd_sc_hd__dfxbp_1 s992 (.CLK(clknet_leaf_28_clk),
    .D(net605),
    .Q(net1085),
    .Q_N(net1084));
 sky130_fd_sc_hd__dfxbp_1 s993 (.CLK(clknet_leaf_31_clk),
    .D(net606),
    .Q(net1087),
    .Q_N(net1086));
 sky130_fd_sc_hd__dfxtp_2 s994 (.CLK(clknet_leaf_31_clk),
    .D(net609),
    .Q(net1088));
 sky130_fd_sc_hd__dfxtp_1 s995 (.CLK(clknet_leaf_31_clk),
    .D(net611),
    .Q(net1089));
 sky130_fd_sc_hd__dfxtp_2 s996 (.CLK(clknet_leaf_27_clk),
    .D(net613),
    .Q(net1090));
 sky130_fd_sc_hd__dlclkp_1 s997 (.CLK(clknet_leaf_26_clk),
    .GATE(net614),
    .GCLK(net1091));
 sky130_fd_sc_hd__dlclkp_2 s998 (.CLK(clknet_leaf_33_clk),
    .GATE(net629),
    .GCLK(net1092));
 sky130_fd_sc_hd__dlclkp_4 s999 (.CLK(clknet_leaf_33_clk),
    .GATE(net634),
    .GCLK(net1093));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(in0),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(in1),
    .X(net754));
 sky130_fd_sc_hd__buf_1 input3 (.A(in10),
    .X(net765));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(in11),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(in12),
    .X(net781));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(in13),
    .X(net794));
 sky130_fd_sc_hd__buf_1 input7 (.A(in14),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(in15),
    .X(net1129));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(in16),
    .X(net1130));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(in17),
    .X(net1131));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(in18),
    .X(net1132));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(in19),
    .X(net1133));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(in2),
    .X(net1134));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(in20),
    .X(net1135));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(in21),
    .X(net1136));
 sky130_fd_sc_hd__buf_1 input16 (.A(in22),
    .X(net1137));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(in23),
    .X(net1138));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(in24),
    .X(net1139));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(in3),
    .X(net1140));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(in4),
    .X(net1141));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(in5),
    .X(net1142));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(in6),
    .X(net1143));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(in7),
    .X(net1144));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(in8),
    .X(net1145));
 sky130_fd_sc_hd__buf_1 input25 (.A(in9),
    .X(net1146));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net1147),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output27 (.A(net1148),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output28 (.A(net1149),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(clknet_1_0__leaf_net1150),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output30 (.A(net1151),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output31 (.A(net1152),
    .X(out14));
 sky130_fd_sc_hd__clkbuf_1 output32 (.A(clknet_1_1__leaf_net1153),
    .X(out15));
 sky130_fd_sc_hd__buf_8 output33 (.A(clknet_1_0__leaf_net1154),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output34 (.A(net1155),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output35 (.A(net1156),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output36 (.A(net1157),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output37 (.A(net1158),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output38 (.A(net1159),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_1 output39 (.A(clknet_1_1__leaf_net1160),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output40 (.A(net1161),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output41 (.A(net1185),
    .X(out9));
 sky130_fd_sc_hd__buf_2 fanout42 (.A(net464),
    .X(net1163));
 sky130_fd_sc_hd__clkbuf_2 fanout43 (.A(net374),
    .X(net1164));
 sky130_fd_sc_hd__buf_2 fanout44 (.A(net271),
    .X(net1165));
 sky130_fd_sc_hd__buf_2 fanout45 (.A(net21),
    .X(net1166));
 sky130_fd_sc_hd__clkbuf_2 fanout46 (.A(net1168),
    .X(net1167));
 sky130_fd_sc_hd__clkbuf_2 fanout47 (.A(net201),
    .X(net1168));
 sky130_fd_sc_hd__clkbuf_2 fanout48 (.A(net1170),
    .X(net1169));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout49 (.A(net1171),
    .X(net1170));
 sky130_fd_sc_hd__clkbuf_2 fanout50 (.A(net62),
    .X(net1171));
 sky130_fd_sc_hd__clkbuf_2 fanout51 (.A(net1173),
    .X(net1172));
 sky130_fd_sc_hd__buf_2 fanout52 (.A(net578),
    .X(net1173));
 sky130_fd_sc_hd__clkbuf_2 fanout53 (.A(net20),
    .X(net1174));
 sky130_fd_sc_hd__buf_2 fanout54 (.A(net372),
    .X(net1175));
 sky130_fd_sc_hd__buf_2 fanout55 (.A(net1177),
    .X(net1176));
 sky130_fd_sc_hd__buf_2 fanout56 (.A(net323),
    .X(net1177));
 sky130_fd_sc_hd__buf_2 fanout57 (.A(net274),
    .X(net1178));
 sky130_fd_sc_hd__buf_2 fanout58 (.A(net89),
    .X(net1179));
 sky130_fd_sc_hd__clkbuf_2 fanout59 (.A(net42),
    .X(net1180));
 sky130_fd_sc_hd__buf_2 fanout60 (.A(net644),
    .X(net1181));
 sky130_fd_sc_hd__buf_2 fanout61 (.A(net1183),
    .X(net1182));
 sky130_fd_sc_hd__clkbuf_2 fanout62 (.A(net643),
    .X(net1183));
 sky130_fd_sc_hd__clkbuf_2 fanout63 (.A(net620),
    .X(net1184));
 sky130_fd_sc_hd__clkbuf_2 fanout64 (.A(net1162),
    .X(net1185));
 sky130_fd_sc_hd__clkbuf_2 fanout65 (.A(net441),
    .X(net1186));
 sky130_fd_sc_hd__buf_1 fanout66 (.A(net441),
    .X(net1187));
 sky130_fd_sc_hd__clkbuf_2 fanout67 (.A(net440),
    .X(net1188));
 sky130_fd_sc_hd__buf_1 fanout68 (.A(net440),
    .X(net1189));
 sky130_fd_sc_hd__buf_2 fanout69 (.A(net421),
    .X(net1190));
 sky130_fd_sc_hd__clkbuf_4 fanout70 (.A(net1192),
    .X(net1191));
 sky130_fd_sc_hd__clkbuf_2 fanout71 (.A(net397),
    .X(net1192));
 sky130_fd_sc_hd__clkbuf_2 fanout72 (.A(net1194),
    .X(net1193));
 sky130_fd_sc_hd__clkbuf_2 fanout73 (.A(net1195),
    .X(net1194));
 sky130_fd_sc_hd__clkbuf_2 fanout74 (.A(net293),
    .X(net1195));
 sky130_fd_sc_hd__buf_2 max_cap75 (.A(net1215),
    .X(net1196));
 sky130_fd_sc_hd__buf_2 fanout76 (.A(net1042),
    .X(net1197));
 sky130_fd_sc_hd__buf_2 fanout77 (.A(net1029),
    .X(net1198));
 sky130_fd_sc_hd__clkbuf_4 fanout78 (.A(net1000),
    .X(net1199));
 sky130_fd_sc_hd__clkbuf_4 fanout79 (.A(net987),
    .X(net1200));
 sky130_fd_sc_hd__clkbuf_4 fanout80 (.A(net986),
    .X(net1201));
 sky130_fd_sc_hd__clkbuf_4 fanout81 (.A(net1277),
    .X(net1202));
 sky130_fd_sc_hd__buf_2 fanout82 (.A(net903),
    .X(net1203));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout83 (.A(net903),
    .X(net1204));
 sky130_fd_sc_hd__clkbuf_4 fanout84 (.A(net1098),
    .X(net1205));
 sky130_fd_sc_hd__clkbuf_2 fanout85 (.A(net731),
    .X(net1206));
 sky130_fd_sc_hd__clkbuf_2 fanout86 (.A(net107),
    .X(net1207));
 sky130_fd_sc_hd__buf_1 fanout87 (.A(net107),
    .X(net1208));
 sky130_fd_sc_hd__clkbuf_4 fanout88 (.A(net742),
    .X(net1209));
 sky130_fd_sc_hd__buf_2 fanout89 (.A(net396),
    .X(net1210));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_36_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_37_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_38_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_39_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_40_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_41_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_42_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_43_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_44_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_45_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_46_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_47_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_48_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1093 (.A(net1093),
    .X(clknet_0_net1093));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1093 (.A(clknet_0_net1093),
    .X(clknet_1_0__leaf_net1093));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1093 (.A(clknet_0_net1093),
    .X(clknet_1_1__leaf_net1093));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1154 (.A(net1154),
    .X(clknet_0_net1154));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1154 (.A(clknet_0_net1154),
    .X(clknet_1_0__leaf_net1154));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1154 (.A(clknet_0_net1154),
    .X(clknet_1_1__leaf_net1154));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1092 (.A(net1092),
    .X(clknet_0_net1092));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1092 (.A(clknet_0_net1092),
    .X(clknet_1_0__leaf_net1092));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1092 (.A(clknet_0_net1092),
    .X(clknet_1_1__leaf_net1092));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net886 (.A(net886),
    .X(clknet_0_net886));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net886 (.A(clknet_0_net886),
    .X(clknet_1_0__leaf_net886));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net886 (.A(clknet_0_net886),
    .X(clknet_1_1__leaf_net886));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1091 (.A(net1091),
    .X(clknet_0_net1091));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1091 (.A(clknet_0_net1091),
    .X(clknet_1_0__leaf_net1091));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1091 (.A(clknet_0_net1091),
    .X(clknet_1_1__leaf_net1091));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net848 (.A(net848),
    .X(clknet_0_net848));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net848 (.A(clknet_0_net848),
    .X(clknet_1_0__leaf_net848));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net848 (.A(clknet_0_net848),
    .X(clknet_1_1__leaf_net848));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net608 (.A(net608),
    .X(clknet_0_net608));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net608 (.A(clknet_0_net608),
    .X(clknet_1_0__leaf_net608));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net608 (.A(clknet_0_net608),
    .X(clknet_1_1__leaf_net608));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net615 (.A(net615),
    .X(clknet_0_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net615 (.A(clknet_0_net615),
    .X(clknet_1_0__leaf_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net615 (.A(clknet_0_net615),
    .X(clknet_1_1__leaf_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net892 (.A(net892),
    .X(clknet_0_net892));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net892 (.A(clknet_0_net892),
    .X(clknet_1_0__leaf_net892));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net892 (.A(clknet_0_net892),
    .X(clknet_1_1__leaf_net892));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1153 (.A(net1153),
    .X(clknet_0_net1153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1153 (.A(clknet_0_net1153),
    .X(clknet_1_0__leaf_net1153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1153 (.A(clknet_0_net1153),
    .X(clknet_1_1__leaf_net1153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net507 (.A(net507),
    .X(clknet_0_net507));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net507 (.A(clknet_0_net507),
    .X(clknet_1_0__leaf_net507));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net507 (.A(clknet_0_net507),
    .X(clknet_1_1__leaf_net507));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1160 (.A(net1160),
    .X(clknet_0_net1160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1160 (.A(clknet_0_net1160),
    .X(clknet_1_0__leaf_net1160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1160 (.A(clknet_0_net1160),
    .X(clknet_1_1__leaf_net1160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1150 (.A(net1150),
    .X(clknet_0_net1150));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1150 (.A(clknet_0_net1150),
    .X(clknet_1_0__leaf_net1150));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1150 (.A(clknet_0_net1150),
    .X(clknet_1_1__leaf_net1150));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1072 (.A(net1072),
    .X(clknet_0_net1072));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1072 (.A(clknet_0_net1072),
    .X(clknet_1_0__leaf_net1072));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1072 (.A(clknet_0_net1072),
    .X(clknet_1_1__leaf_net1072));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net574 (.A(net574),
    .X(clknet_0_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net574 (.A(clknet_0_net574),
    .X(clknet_1_0__leaf_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net574 (.A(clknet_0_net574),
    .X(clknet_1_1__leaf_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1109 (.A(net1109),
    .X(clknet_0_net1109));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1109 (.A(clknet_0_net1109),
    .X(clknet_1_0__leaf_net1109));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1109 (.A(clknet_0_net1109),
    .X(clknet_1_1__leaf_net1109));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1111 (.A(net1111),
    .X(clknet_0_net1111));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1111 (.A(clknet_0_net1111),
    .X(clknet_1_0__leaf_net1111));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1111 (.A(clknet_0_net1111),
    .X(clknet_1_1__leaf_net1111));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net689 (.A(net689),
    .X(clknet_0_net689));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net689 (.A(clknet_0_net689),
    .X(clknet_1_0__leaf_net689));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net689 (.A(clknet_0_net689),
    .X(clknet_1_1__leaf_net689));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net570 (.A(net570),
    .X(clknet_0_net570));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net570 (.A(clknet_0_net570),
    .X(clknet_1_0__leaf_net570));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net570 (.A(clknet_0_net570),
    .X(clknet_1_1__leaf_net570));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1071 (.A(net1071),
    .X(clknet_0_net1071));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1071 (.A(clknet_0_net1071),
    .X(clknet_1_0__leaf_net1071));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1071 (.A(clknet_0_net1071),
    .X(clknet_1_1__leaf_net1071));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1070 (.A(net1070),
    .X(clknet_0_net1070));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1070 (.A(clknet_0_net1070),
    .X(clknet_1_0__leaf_net1070));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1070 (.A(clknet_0_net1070),
    .X(clknet_1_1__leaf_net1070));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1052 (.A(net1052),
    .X(clknet_0_net1052));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1052 (.A(clknet_0_net1052),
    .X(clknet_1_0__leaf_net1052));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1052 (.A(clknet_0_net1052),
    .X(clknet_1_1__leaf_net1052));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1051 (.A(net1051),
    .X(clknet_0_net1051));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1051 (.A(clknet_0_net1051),
    .X(clknet_1_0__leaf_net1051));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1051 (.A(clknet_0_net1051),
    .X(clknet_1_1__leaf_net1051));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1050 (.A(net1050),
    .X(clknet_0_net1050));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1050 (.A(clknet_0_net1050),
    .X(clknet_1_0__leaf_net1050));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1050 (.A(clknet_0_net1050),
    .X(clknet_1_1__leaf_net1050));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net524 (.A(net524),
    .X(clknet_0_net524));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net524 (.A(clknet_0_net524),
    .X(clknet_1_0__leaf_net524));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net524 (.A(clknet_0_net524),
    .X(clknet_1_1__leaf_net524));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1032 (.A(net1032),
    .X(clknet_0_net1032));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1032 (.A(clknet_0_net1032),
    .X(clknet_1_0__leaf_net1032));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1032 (.A(clknet_0_net1032),
    .X(clknet_1_1__leaf_net1032));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net458 (.A(net458),
    .X(clknet_0_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net458 (.A(clknet_0_net458),
    .X(clknet_1_0__leaf_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net458 (.A(clknet_0_net458),
    .X(clknet_1_1__leaf_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1031 (.A(net1031),
    .X(clknet_0_net1031));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1031 (.A(clknet_0_net1031),
    .X(clknet_1_0__leaf_net1031));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1031 (.A(clknet_0_net1031),
    .X(clknet_1_1__leaf_net1031));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net457 (.A(net457),
    .X(clknet_0_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net457 (.A(clknet_0_net457),
    .X(clknet_1_0__leaf_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net457 (.A(clknet_0_net457),
    .X(clknet_1_1__leaf_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1030 (.A(net1030),
    .X(clknet_0_net1030));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1030 (.A(clknet_0_net1030),
    .X(clknet_1_0__leaf_net1030));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1030 (.A(clknet_0_net1030),
    .X(clknet_1_1__leaf_net1030));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1011 (.A(net1011),
    .X(clknet_0_net1011));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1011 (.A(clknet_0_net1011),
    .X(clknet_1_0__leaf_net1011));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1011 (.A(clknet_0_net1011),
    .X(clknet_1_1__leaf_net1011));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1010 (.A(net1010),
    .X(clknet_0_net1010));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1010 (.A(clknet_0_net1010),
    .X(clknet_1_0__leaf_net1010));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1010 (.A(clknet_0_net1010),
    .X(clknet_1_1__leaf_net1010));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net381 (.A(net381),
    .X(clknet_0_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net381 (.A(clknet_0_net381),
    .X(clknet_1_0__leaf_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net381 (.A(clknet_0_net381),
    .X(clknet_1_1__leaf_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net385 (.A(net385),
    .X(clknet_0_net385));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net385 (.A(clknet_0_net385),
    .X(clknet_1_0__leaf_net385));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net385 (.A(clknet_0_net385),
    .X(clknet_1_1__leaf_net385));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1009 (.A(net1009),
    .X(clknet_0_net1009));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1009 (.A(clknet_0_net1009),
    .X(clknet_1_0__leaf_net1009));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1009 (.A(clknet_0_net1009),
    .X(clknet_1_1__leaf_net1009));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net990 (.A(net990),
    .X(clknet_0_net990));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net990 (.A(clknet_0_net990),
    .X(clknet_1_0__leaf_net990));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net990 (.A(clknet_0_net990),
    .X(clknet_1_1__leaf_net990));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net417 (.A(net417),
    .X(clknet_0_net417));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net417 (.A(clknet_0_net417),
    .X(clknet_1_0__leaf_net417));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net417 (.A(clknet_0_net417),
    .X(clknet_1_1__leaf_net417));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net418 (.A(net418),
    .X(clknet_0_net418));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net418 (.A(clknet_0_net418),
    .X(clknet_1_0__leaf_net418));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net418 (.A(clknet_0_net418),
    .X(clknet_1_1__leaf_net418));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net290 (.A(net290),
    .X(clknet_0_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net290 (.A(clknet_0_net290),
    .X(clknet_1_0__leaf_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net290 (.A(clknet_0_net290),
    .X(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net989 (.A(net989),
    .X(clknet_0_net989));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net989 (.A(clknet_0_net989),
    .X(clknet_1_0__leaf_net989));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net989 (.A(clknet_0_net989),
    .X(clknet_1_1__leaf_net989));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net988 (.A(net988),
    .X(clknet_0_net988));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net988 (.A(clknet_0_net988),
    .X(clknet_1_0__leaf_net988));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net988 (.A(clknet_0_net988),
    .X(clknet_1_1__leaf_net988));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net969 (.A(net969),
    .X(clknet_0_net969));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net969 (.A(clknet_0_net969),
    .X(clknet_1_0__leaf_net969));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net969 (.A(clknet_0_net969),
    .X(clknet_1_1__leaf_net969));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net341 (.A(net341),
    .X(clknet_0_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net341 (.A(clknet_0_net341),
    .X(clknet_1_0__leaf_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net341 (.A(clknet_0_net341),
    .X(clknet_1_1__leaf_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net228 (.A(net228),
    .X(clknet_0_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net228 (.A(clknet_0_net228),
    .X(clknet_1_0__leaf_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net228 (.A(clknet_0_net228),
    .X(clknet_1_1__leaf_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net968 (.A(net968),
    .X(clknet_0_net968));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net968 (.A(clknet_0_net968),
    .X(clknet_1_0__leaf_net968));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net968 (.A(clknet_0_net968),
    .X(clknet_1_1__leaf_net968));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net487 (.A(net487),
    .X(clknet_0_net487));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net487 (.A(clknet_0_net487),
    .X(clknet_1_0__leaf_net487));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net487 (.A(clknet_0_net487),
    .X(clknet_1_1__leaf_net487));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net503 (.A(net503),
    .X(clknet_0_net503));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net503 (.A(clknet_0_net503),
    .X(clknet_1_0__leaf_net503));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net503 (.A(clknet_0_net503),
    .X(clknet_1_1__leaf_net503));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net499 (.A(net499),
    .X(clknet_0_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net499 (.A(clknet_0_net499),
    .X(clknet_1_0__leaf_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net499 (.A(clknet_0_net499),
    .X(clknet_1_1__leaf_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net492 (.A(net492),
    .X(clknet_0_net492));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net492 (.A(clknet_0_net492),
    .X(clknet_1_0__leaf_net492));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net492 (.A(clknet_0_net492),
    .X(clknet_1_1__leaf_net492));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net489 (.A(net489),
    .X(clknet_0_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_0__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_1__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net488 (.A(net488),
    .X(clknet_0_net488));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net488 (.A(clknet_0_net488),
    .X(clknet_1_0__leaf_net488));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net488 (.A(clknet_0_net488),
    .X(clknet_1_1__leaf_net488));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net238 (.A(net238),
    .X(clknet_0_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net238 (.A(clknet_0_net238),
    .X(clknet_1_0__leaf_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net238 (.A(clknet_0_net238),
    .X(clknet_1_1__leaf_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net227 (.A(net227),
    .X(clknet_0_net227));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net227 (.A(clknet_0_net227),
    .X(clknet_1_0__leaf_net227));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net227 (.A(clknet_0_net227),
    .X(clknet_1_1__leaf_net227));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net226 (.A(net226),
    .X(clknet_0_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net226 (.A(clknet_0_net226),
    .X(clknet_1_0__leaf_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net226 (.A(clknet_0_net226),
    .X(clknet_1_1__leaf_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net967 (.A(net967),
    .X(clknet_0_net967));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net967 (.A(clknet_0_net967),
    .X(clknet_1_0__leaf_net967));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net967 (.A(clknet_0_net967),
    .X(clknet_1_1__leaf_net967));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net948 (.A(net948),
    .X(clknet_0_net948));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net948 (.A(clknet_0_net948),
    .X(clknet_1_0__leaf_net948));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net948 (.A(clknet_0_net948),
    .X(clknet_1_1__leaf_net948));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net297 (.A(net297),
    .X(clknet_0_net297));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net297 (.A(clknet_0_net297),
    .X(clknet_1_0__leaf_net297));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net297 (.A(clknet_0_net297),
    .X(clknet_1_1__leaf_net297));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net891 (.A(net891),
    .X(clknet_0_net891));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net891 (.A(clknet_0_net891),
    .X(clknet_1_0__leaf_net891));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net891 (.A(clknet_0_net891),
    .X(clknet_1_1__leaf_net891));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net595 (.A(net595),
    .X(clknet_0_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net595 (.A(net1211),
    .X(clknet_1_0__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_1__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net692 (.A(net692),
    .X(clknet_0_net692));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net692 (.A(clknet_0_net692),
    .X(clknet_1_0__leaf_net692));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net692 (.A(clknet_0_net692),
    .X(clknet_1_1__leaf_net692));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net694 (.A(net694),
    .X(clknet_0_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net694 (.A(clknet_0_net694),
    .X(clknet_1_0__leaf_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net694 (.A(clknet_0_net694),
    .X(clknet_1_1__leaf_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net618 (.A(net618),
    .X(clknet_0_net618));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net618 (.A(clknet_0_net618),
    .X(clknet_1_0__leaf_net618));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net618 (.A(net1213),
    .X(clknet_1_1__leaf_net618));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net619 (.A(net619),
    .X(clknet_0_net619));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net619 (.A(clknet_0_net619),
    .X(clknet_1_0__leaf_net619));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net619 (.A(clknet_0_net619),
    .X(clknet_1_1__leaf_net619));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net596 (.A(net596),
    .X(clknet_0_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net596 (.A(clknet_0_net596),
    .X(clknet_1_0__leaf_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net596 (.A(clknet_0_net596),
    .X(clknet_1_1__leaf_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net202 (.A(net202),
    .X(clknet_0_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net202 (.A(clknet_0_net202),
    .X(clknet_1_0__leaf_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net202 (.A(clknet_0_net202),
    .X(clknet_1_1__leaf_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net220 (.A(net220),
    .X(clknet_0_net220));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net220 (.A(clknet_0_net220),
    .X(clknet_1_0__leaf_net220));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net220 (.A(clknet_0_net220),
    .X(clknet_1_1__leaf_net220));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net846 (.A(net846),
    .X(clknet_0_net846));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net846 (.A(clknet_0_net846),
    .X(clknet_1_0__leaf_net846));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net846 (.A(clknet_0_net846),
    .X(clknet_1_1__leaf_net846));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net216 (.A(net216),
    .X(clknet_0_net216));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net216 (.A(clknet_0_net216),
    .X(clknet_1_0__leaf_net216));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net216 (.A(clknet_0_net216),
    .X(clknet_1_1__leaf_net216));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net211 (.A(net211),
    .X(clknet_0_net211));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net211 (.A(clknet_0_net211),
    .X(clknet_1_0__leaf_net211));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net211 (.A(clknet_0_net211),
    .X(clknet_1_1__leaf_net211));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net210 (.A(net210),
    .X(clknet_0_net210));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net210 (.A(clknet_0_net210),
    .X(clknet_1_0__leaf_net210));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net210 (.A(clknet_0_net210),
    .X(clknet_1_1__leaf_net210));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net208 (.A(net208),
    .X(clknet_0_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net208 (.A(clknet_0_net208),
    .X(clknet_1_0__leaf_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net208 (.A(clknet_0_net208),
    .X(clknet_1_1__leaf_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net205 (.A(net205),
    .X(clknet_0_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net205 (.A(clknet_0_net205),
    .X(clknet_1_0__leaf_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net205 (.A(clknet_0_net205),
    .X(clknet_1_1__leaf_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net204 (.A(net204),
    .X(clknet_0_net204));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net204 (.A(clknet_0_net204),
    .X(clknet_1_0__leaf_net204));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net204 (.A(clknet_0_net204),
    .X(clknet_1_1__leaf_net204));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net203 (.A(net203),
    .X(clknet_0_net203));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net203 (.A(clknet_0_net203),
    .X(clknet_1_0__leaf_net203));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net203 (.A(clknet_0_net203),
    .X(clknet_1_1__leaf_net203));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net298 (.A(net298),
    .X(clknet_0_net298));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net298 (.A(clknet_0_net298),
    .X(clknet_1_0__leaf_net298));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net298 (.A(clknet_0_net298),
    .X(clknet_1_1__leaf_net298));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net890 (.A(net890),
    .X(clknet_0_net890));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net890 (.A(clknet_0_net890),
    .X(clknet_1_0__leaf_net890));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net890 (.A(clknet_0_net890),
    .X(clknet_1_1__leaf_net890));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net469 (.A(net469),
    .X(clknet_0_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net469 (.A(clknet_0_net469),
    .X(clknet_1_0__leaf_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net469 (.A(clknet_0_net469),
    .X(clknet_1_1__leaf_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net483 (.A(net483),
    .X(clknet_0_net483));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net483 (.A(clknet_0_net483),
    .X(clknet_1_0__leaf_net483));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net483 (.A(clknet_0_net483),
    .X(clknet_1_1__leaf_net483));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net479 (.A(net479),
    .X(clknet_0_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net479 (.A(clknet_0_net479),
    .X(clknet_1_0__leaf_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net479 (.A(clknet_0_net479),
    .X(clknet_1_1__leaf_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net482 (.A(net482),
    .X(clknet_0_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net482 (.A(clknet_0_net482),
    .X(clknet_1_0__leaf_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net482 (.A(clknet_0_net482),
    .X(clknet_1_1__leaf_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net465 (.A(net465),
    .X(clknet_0_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net465 (.A(clknet_0_net465),
    .X(clknet_1_0__leaf_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net465 (.A(clknet_0_net465),
    .X(clknet_1_1__leaf_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net947 (.A(net947),
    .X(clknet_0_net947));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net947 (.A(clknet_0_net947),
    .X(clknet_1_0__leaf_net947));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net947 (.A(clknet_0_net947),
    .X(clknet_1_1__leaf_net947));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net200 (.A(net200),
    .X(clknet_0_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net200 (.A(clknet_0_net200),
    .X(clknet_1_0__leaf_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net200 (.A(clknet_0_net200),
    .X(clknet_1_1__leaf_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net318 (.A(net318),
    .X(clknet_0_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net318 (.A(clknet_0_net318),
    .X(clknet_1_0__leaf_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net318 (.A(clknet_0_net318),
    .X(clknet_1_1__leaf_net318));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net180 (.A(net180),
    .X(clknet_0_net180));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net180 (.A(clknet_0_net180),
    .X(clknet_1_0__leaf_net180));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net180 (.A(clknet_0_net180),
    .X(clknet_1_1__leaf_net180));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net195 (.A(net195),
    .X(clknet_0_net195));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net195 (.A(clknet_0_net195),
    .X(clknet_1_0__leaf_net195));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net195 (.A(clknet_0_net195),
    .X(clknet_1_1__leaf_net195));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net185 (.A(net185),
    .X(clknet_0_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net185 (.A(clknet_0_net185),
    .X(clknet_1_0__leaf_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net185 (.A(clknet_0_net185),
    .X(clknet_1_1__leaf_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net181 (.A(net181),
    .X(clknet_0_net181));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net181 (.A(clknet_0_net181),
    .X(clknet_1_0__leaf_net181));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net181 (.A(clknet_0_net181),
    .X(clknet_1_1__leaf_net181));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net179 (.A(net179),
    .X(clknet_0_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_0__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_1__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net946 (.A(net946),
    .X(clknet_0_net946));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net946 (.A(clknet_0_net946),
    .X(clknet_1_0__leaf_net946));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net946 (.A(clknet_0_net946),
    .X(clknet_1_1__leaf_net946));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net927 (.A(net927),
    .X(clknet_0_net927));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net927 (.A(clknet_0_net927),
    .X(clknet_1_0__leaf_net927));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net927 (.A(clknet_0_net927),
    .X(clknet_1_1__leaf_net927));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net248 (.A(net248),
    .X(clknet_0_net248));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net248 (.A(clknet_0_net248),
    .X(clknet_1_0__leaf_net248));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net248 (.A(clknet_0_net248),
    .X(clknet_1_1__leaf_net248));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net260 (.A(net260),
    .X(clknet_0_net260));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net260 (.A(clknet_0_net260),
    .X(clknet_1_0__leaf_net260));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net260 (.A(clknet_0_net260),
    .X(clknet_1_1__leaf_net260));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net252 (.A(net252),
    .X(clknet_0_net252));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net252 (.A(clknet_0_net252),
    .X(clknet_1_0__leaf_net252));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net252 (.A(clknet_0_net252),
    .X(clknet_1_1__leaf_net252));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net249 (.A(net249),
    .X(clknet_0_net249));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net249 (.A(clknet_0_net249),
    .X(clknet_1_0__leaf_net249));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net249 (.A(clknet_0_net249),
    .X(clknet_1_1__leaf_net249));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net247 (.A(net247),
    .X(clknet_0_net247));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net247 (.A(clknet_0_net247),
    .X(clknet_1_0__leaf_net247));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net247 (.A(clknet_0_net247),
    .X(clknet_1_1__leaf_net247));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net127 (.A(net127),
    .X(clknet_0_net127));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net127 (.A(clknet_0_net127),
    .X(clknet_1_0__leaf_net127));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net127 (.A(clknet_0_net127),
    .X(clknet_1_1__leaf_net127));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net926 (.A(net926),
    .X(clknet_0_net926));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net926 (.A(clknet_0_net926),
    .X(clknet_1_0__leaf_net926));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net926 (.A(clknet_0_net926),
    .X(clknet_1_1__leaf_net926));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net925 (.A(net925),
    .X(clknet_0_net925));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net925 (.A(clknet_0_net925),
    .X(clknet_1_0__leaf_net925));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net925 (.A(clknet_0_net925),
    .X(clknet_1_1__leaf_net925));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net105 (.A(net105),
    .X(clknet_0_net105));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net105 (.A(clknet_0_net105),
    .X(clknet_1_0__leaf_net105));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net105 (.A(clknet_0_net105),
    .X(clknet_1_1__leaf_net105));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net906 (.A(net906),
    .X(clknet_0_net906));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net906 (.A(clknet_0_net906),
    .X(clknet_1_0__leaf_net906));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net906 (.A(clknet_0_net906),
    .X(clknet_1_1__leaf_net906));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net37 (.A(net37),
    .X(clknet_0_net37));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net37 (.A(clknet_0_net37),
    .X(clknet_1_0__leaf_net37));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net37 (.A(clknet_0_net37),
    .X(clknet_1_1__leaf_net37));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net35 (.A(net35),
    .X(clknet_0_net35));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net35 (.A(clknet_0_net35),
    .X(clknet_1_0__leaf_net35));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net35 (.A(clknet_0_net35),
    .X(clknet_1_1__leaf_net35));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net905 (.A(net905),
    .X(clknet_0_net905));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net905 (.A(clknet_0_net905),
    .X(clknet_1_0__leaf_net905));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net905 (.A(clknet_0_net905),
    .X(clknet_1_1__leaf_net905));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net157 (.A(net157),
    .X(clknet_0_net157));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net157 (.A(clknet_0_net157),
    .X(clknet_1_0__leaf_net157));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net157 (.A(clknet_0_net157),
    .X(clknet_1_1__leaf_net157));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net155 (.A(net155),
    .X(clknet_0_net155));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net155 (.A(clknet_0_net155),
    .X(clknet_1_0__leaf_net155));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net155 (.A(clknet_0_net155),
    .X(clknet_1_1__leaf_net155));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net171 (.A(net171),
    .X(clknet_0_net171));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net171 (.A(clknet_0_net171),
    .X(clknet_1_0__leaf_net171));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net171 (.A(clknet_0_net171),
    .X(clknet_1_1__leaf_net171));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net159 (.A(net159),
    .X(clknet_0_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net159 (.A(clknet_0_net159),
    .X(clknet_1_0__leaf_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net159 (.A(clknet_0_net159),
    .X(clknet_1_1__leaf_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net156 (.A(net156),
    .X(clknet_0_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net156 (.A(clknet_0_net156),
    .X(clknet_1_0__leaf_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net156 (.A(clknet_0_net156),
    .X(clknet_1_1__leaf_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net904 (.A(net904),
    .X(clknet_0_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net904 (.A(clknet_0_net904),
    .X(clknet_1_0__leaf_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net904 (.A(clknet_0_net904),
    .X(clknet_1_1__leaf_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1128 (.A(net1128),
    .X(clknet_0_net1128));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1128 (.A(clknet_0_net1128),
    .X(clknet_1_0__leaf_net1128));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1128 (.A(clknet_0_net1128),
    .X(clknet_1_1__leaf_net1128));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net533 (.A(net533),
    .X(clknet_0_net533));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net533 (.A(clknet_0_net533),
    .X(clknet_1_0__leaf_net533));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net533 (.A(clknet_0_net533),
    .X(clknet_1_1__leaf_net533));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net548 (.A(net548),
    .X(clknet_0_net548));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net548 (.A(clknet_0_net548),
    .X(clknet_1_0__leaf_net548));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net548 (.A(clknet_0_net548),
    .X(clknet_1_1__leaf_net548));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net667 (.A(net667),
    .X(clknet_0_net667));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net667 (.A(clknet_0_net667),
    .X(clknet_1_0__leaf_net667));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net667 (.A(clknet_0_net667),
    .X(clknet_1_1__leaf_net667));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net681 (.A(net681),
    .X(clknet_0_net681));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net681 (.A(clknet_0_net681),
    .X(clknet_1_0__leaf_net681));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net681 (.A(clknet_0_net681),
    .X(clknet_1_1__leaf_net681));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1110 (.A(net1110),
    .X(clknet_0_net1110));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1110 (.A(clknet_0_net1110),
    .X(clknet_1_0__leaf_net1110));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1110 (.A(clknet_0_net1110),
    .X(clknet_1_1__leaf_net1110));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net668 (.A(net668),
    .X(clknet_0_net668));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net668 (.A(clknet_0_net668),
    .X(clknet_1_0__leaf_net668));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net668 (.A(clknet_0_net668),
    .X(clknet_1_1__leaf_net668));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net641 (.A(net641),
    .X(clknet_0_net641));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net641 (.A(clknet_0_net641),
    .X(clknet_1_0__leaf_net641));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net641 (.A(clknet_0_net641),
    .X(clknet_1_1__leaf_net641));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net642 (.A(net642),
    .X(clknet_0_net642));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net642 (.A(clknet_0_net642),
    .X(clknet_1_0__leaf_net642));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net642 (.A(clknet_0_net642),
    .X(clknet_1_1__leaf_net642));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net553 (.A(net553),
    .X(clknet_0_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net553 (.A(clknet_0_net553),
    .X(clknet_1_0__leaf_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net553 (.A(clknet_0_net553),
    .X(clknet_1_1__leaf_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net554 (.A(net554),
    .X(clknet_0_net554));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net554 (.A(clknet_0_net554),
    .X(clknet_1_0__leaf_net554));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net554 (.A(clknet_0_net554),
    .X(clknet_1_1__leaf_net554));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net549 (.A(net549),
    .X(clknet_0_net549));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net549 (.A(clknet_0_net549),
    .X(clknet_1_0__leaf_net549));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net549 (.A(clknet_0_net549),
    .X(clknet_1_1__leaf_net549));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net550 (.A(net550),
    .X(clknet_0_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net550 (.A(clknet_0_net550),
    .X(clknet_1_0__leaf_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net550 (.A(clknet_0_net550),
    .X(clknet_1_1__leaf_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net535 (.A(net535),
    .X(clknet_0_net535));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net535 (.A(clknet_0_net535),
    .X(clknet_1_0__leaf_net535));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net535 (.A(clknet_0_net535),
    .X(clknet_1_1__leaf_net535));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net539 (.A(net539),
    .X(clknet_0_net539));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net539 (.A(clknet_0_net539),
    .X(clknet_1_0__leaf_net539));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net539 (.A(clknet_0_net539),
    .X(clknet_1_1__leaf_net539));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net278 (.A(net278),
    .X(clknet_0_net278));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net278 (.A(clknet_0_net278),
    .X(clknet_1_0__leaf_net278));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net278 (.A(clknet_0_net278),
    .X(clknet_1_1__leaf_net278));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net855 (.A(net855),
    .X(clknet_0_net855));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net855 (.A(clknet_0_net855),
    .X(clknet_1_0__leaf_net855));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net855 (.A(clknet_0_net855),
    .X(clknet_1_1__leaf_net855));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(clknet_0_net595),
    .X(net1211));
 sky130_fd_sc_hd__clkbuf_1 clone2 (.A(clknet_0_net618),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(clknet_0_net618),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(clknet_1_1__leaf_net595),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net1061),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net225),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net158),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net224),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net739),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net398),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net713),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net726),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net1007),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net366),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net982),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net817),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net558),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net715),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net993),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net371),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net1090),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net723),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net1115),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net1097),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net1203),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net303),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net394),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net1080),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net991),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net1020),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net1056),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net1035),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net93),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net985),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net136),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net994),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net987),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net343),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net556),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net322),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net1039),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net651),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net138),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net467),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net722),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net255),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net937),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net472),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net1081),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net251),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net1022),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net308),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net319),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net351),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net1027),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net986),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net698),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net349),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net620),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net534),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net1005),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net646),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net345),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net934),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net935),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net719),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net980),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net1065),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net466),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net1006),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net1026),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net427),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net1206),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net1117),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net1005),
    .X(net1285));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold32_A (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_s953_Q_N (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge740_D1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_S1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S0 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_SCE (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_s990_Q (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_S1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_S1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A2 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_SET_B (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_S1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_S1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_S1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout47_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_A0 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_X (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_D1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_X (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A0 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_Q (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge759_D_N (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge743_RESET_B (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A3 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_SCD (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_SCD (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_Q_N (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A0 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A0 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_B (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_Q (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout56_A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_C (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A0 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_X (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A0 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_B (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_B (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_SCD (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A0 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_X (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S0 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A0 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_SCE (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_X (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c659_A0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A2 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_Q (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A3 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_D (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_A3 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_A0 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_A3 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_SCE (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_D1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_SET_B (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_X (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A3 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge761_B (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge745_D (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_A0 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_X (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A2 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_C (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A0 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A0 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_X (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_S0 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_X (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_X (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_D (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge762_A3 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A1 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A2 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_C (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_SCE (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_SCE (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_X (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge762_A2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_D (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S0 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A0 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_DE (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_B (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_C1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_X (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_Q (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_C (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_Q_N (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_A (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_Q (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_S1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_S0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_SCE (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_Q_N (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_Q_N (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_S0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_s873_Q (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_S1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_S1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_S1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_output28_A (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_Q (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A3 (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A2 (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout44_X (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A0 (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_D1 (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_SCD (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A2 (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A0 (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A1 (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_S1 (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A0 (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_SCD (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_X (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_SCD (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A3 (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S0 (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A1 (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_RESET_B (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout49_A (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_X (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_C_N (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_A (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_B1 (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A1 (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A2 (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A2 (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_B (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A1 (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A2 (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout56_X (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_S1 (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_SET_B (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_SET_B (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_RESET_B (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_RESET_B (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_SCD (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_B1 (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A3 (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge740_C1 (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout55_A (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout57_X (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A1 (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A1 (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_RESET_B (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_C (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_D (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A1 (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A2 (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_S0 (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A3 (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_RESET_B (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_X (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A2 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_C1 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_B (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_B (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A2 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_A (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap75_X (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c648_S0 (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_B (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S1 (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_D1 (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_B (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_B (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_SET_B (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_X (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A1 (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A3 (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A3 (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_SCD (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_C1 (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A2 (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A2 (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_SET_B (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_C (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S1 (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_X (.DIODE(net1198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_B (.DIODE(net1198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A3 (.DIODE(net1198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net1198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A3 (.DIODE(net1198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_S0 (.DIODE(net1198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_S1 (.DIODE(net1198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_S1 (.DIODE(net1198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_B (.DIODE(net1198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S0 (.DIODE(net1198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_S0 (.DIODE(net1198));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_X (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_S0 (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A3 (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_S0 (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_S0 (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_S1 (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_S1 (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_C (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_B (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S0 (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_S1 (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_X (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_SET_B (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A3 (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A3 (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A3 (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_S0 (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_S0 (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_SET_B (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S1 (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_X (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_S0 (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_S0 (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_S1 (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_S1 (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_C_N (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_B (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_S1 (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S1 (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold25_A (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_X (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_S1 (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_B (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_B (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_B (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_C (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_C (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c45_C (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_X (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_X (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_X (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_X (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A (.DIODE(clknet_1_1__leaf_net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_C (.DIODE(clknet_1_1__leaf_net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_SCD (.DIODE(clknet_1_1__leaf_net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_S0 (.DIODE(clknet_1_1__leaf_net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_D (.DIODE(clknet_1_1__leaf_net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A1 (.DIODE(clknet_1_1__leaf_net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge760_SET_B (.DIODE(clknet_1_1__leaf_net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net156_X (.DIODE(clknet_1_1__leaf_net156));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
