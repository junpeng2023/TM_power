module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net165;
 wire net176;
 wire net703;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net818;
 wire clknet_1_0__leaf_net818;
 wire clknet_1_1__leaf_net818;
 wire clknet_0_net615;
 wire clknet_1_0__leaf_net615;
 wire clknet_1_1__leaf_net615;
 wire clknet_0_net817;
 wire clknet_1_0__leaf_net817;
 wire clknet_1_1__leaf_net817;
 wire clknet_0_net608;
 wire clknet_1_0__leaf_net608;
 wire clknet_1_1__leaf_net608;
 wire clknet_0_net600;
 wire clknet_1_0__leaf_net600;
 wire clknet_1_1__leaf_net600;
 wire clknet_0_net711;
 wire clknet_1_0__leaf_net711;
 wire clknet_1_1__leaf_net711;
 wire clknet_0_net611;
 wire clknet_1_0__leaf_net611;
 wire clknet_1_1__leaf_net611;
 wire clknet_0_net577;
 wire clknet_1_0__leaf_net577;
 wire clknet_1_1__leaf_net577;
 wire clknet_0_net798;
 wire clknet_1_0__leaf_net798;
 wire clknet_1_1__leaf_net798;
 wire clknet_0_net511;
 wire clknet_1_0__leaf_net511;
 wire clknet_1_1__leaf_net511;
 wire clknet_0_net797;
 wire clknet_1_0__leaf_net797;
 wire clknet_1_1__leaf_net797;
 wire clknet_0_net602;
 wire clknet_1_0__leaf_net602;
 wire clknet_1_1__leaf_net602;
 wire clknet_0_net495;
 wire clknet_1_0__leaf_net495;
 wire clknet_1_1__leaf_net495;
 wire clknet_0_net502;
 wire clknet_1_0__leaf_net502;
 wire clknet_1_1__leaf_net502;
 wire clknet_0_net796;
 wire clknet_1_0__leaf_net796;
 wire clknet_1_1__leaf_net796;
 wire clknet_0_net777;
 wire clknet_1_0__leaf_net777;
 wire clknet_1_1__leaf_net777;
 wire clknet_0_net398;
 wire clknet_1_0__leaf_net398;
 wire clknet_1_1__leaf_net398;
 wire clknet_0_net610;
 wire clknet_1_0__leaf_net610;
 wire clknet_1_1__leaf_net610;
 wire clknet_0_net420;
 wire clknet_1_0__leaf_net420;
 wire clknet_1_1__leaf_net420;
 wire clknet_0_net391;
 wire clknet_1_0__leaf_net391;
 wire clknet_1_1__leaf_net391;
 wire clknet_0_net389;
 wire clknet_1_0__leaf_net389;
 wire clknet_1_1__leaf_net389;
 wire clknet_0_net776;
 wire clknet_1_0__leaf_net776;
 wire clknet_1_1__leaf_net776;
 wire clknet_0_net775;
 wire clknet_1_0__leaf_net775;
 wire clknet_1_1__leaf_net775;
 wire clknet_0_net595;
 wire clknet_1_0__leaf_net595;
 wire clknet_1_1__leaf_net595;
 wire clknet_0_net901;
 wire clknet_1_0__leaf_net901;
 wire clknet_1_1__leaf_net901;
 wire clknet_0_net186;
 wire clknet_1_0__leaf_net186;
 wire clknet_1_1__leaf_net186;
 wire clknet_0_net910;
 wire clknet_1_0__leaf_net910;
 wire clknet_1_1__leaf_net910;
 wire clknet_0_net179;
 wire clknet_1_0__leaf_net179;
 wire clknet_1_1__leaf_net179;
 wire clknet_0_net180;
 wire clknet_1_0__leaf_net180;
 wire clknet_1_1__leaf_net180;
 wire clknet_0_net759;
 wire clknet_1_0__leaf_net759;
 wire clknet_1_1__leaf_net759;
 wire clknet_0_net924;
 wire clknet_1_0__leaf_net924;
 wire clknet_1_1__leaf_net924;
 wire clknet_0_net905;
 wire clknet_1_0__leaf_net905;
 wire clknet_1_1__leaf_net905;
 wire clknet_0_net177;
 wire clknet_1_0__leaf_net177;
 wire clknet_1_1__leaf_net177;
 wire clknet_0_net902;
 wire clknet_1_0__leaf_net902;
 wire clknet_1_1__leaf_net902;
 wire clknet_0_net709;
 wire clknet_1_0__leaf_net709;
 wire clknet_1_1__leaf_net709;
 wire clknet_0_net758;
 wire clknet_1_0__leaf_net758;
 wire clknet_1_1__leaf_net758;
 wire clknet_0_net281;
 wire clknet_1_0__leaf_net281;
 wire clknet_1_1__leaf_net281;
 wire clknet_0_net911;
 wire clknet_1_0__leaf_net911;
 wire clknet_1_1__leaf_net911;
 wire clknet_0_net276;
 wire clknet_1_0__leaf_net276;
 wire clknet_1_1__leaf_net276;
 wire clknet_0_net170;
 wire clknet_1_0__leaf_net170;
 wire clknet_1_1__leaf_net170;
 wire clknet_0_net744;
 wire clknet_1_0__leaf_net744;
 wire clknet_1_1__leaf_net744;
 wire clknet_0_net532;
 wire clknet_1_0__leaf_net532;
 wire clknet_1_1__leaf_net532;
 wire clknet_0_net879;
 wire clknet_1_0__leaf_net879;
 wire clknet_1_1__leaf_net879;
 wire clknet_0_net710;
 wire clknet_1_0__leaf_net710;
 wire clknet_1_1__leaf_net710;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;

 sky130_fd_sc_hd__and3_2 c100 (.A(net1001),
    .B(net11),
    .C(net1000),
    .X(net37));
 sky130_fd_sc_hd__a2111o_1 c101 (.A1(net36),
    .A2(net35),
    .B1(net11),
    .C1(net834),
    .D1(net34),
    .X(net38));
 sky130_fd_sc_hd__and3_1 c102 (.A(net37),
    .B(net30),
    .C(net29),
    .X(net39));
 sky130_fd_sc_hd__or4bb_2 c103 (.A(net34),
    .B(net32),
    .C_N(net35),
    .D_N(net972),
    .X(net40));
 sky130_fd_sc_hd__mux4_2 c104 (.A0(net38),
    .A1(net33),
    .A2(net1018),
    .A3(net24),
    .S0(net837),
    .S1(net35),
    .X(net41));
 sky130_fd_sc_hd__a2111o_4 c105 (.A1(net36),
    .A2(net29),
    .B1(net31),
    .C1(net1003),
    .D1(net41),
    .X(net42));
 sky130_fd_sc_hd__mux4_2 c106 (.A0(net31),
    .A1(net38),
    .A2(net42),
    .A3(net8),
    .S0(net951),
    .S1(net41),
    .X(net43));
 sky130_fd_sc_hd__a2111o_4 c107 (.A1(net28),
    .A2(net871),
    .B1(net42),
    .C1(net856),
    .D1(net43),
    .X(net884));
 sky130_fd_sc_hd__mux4_2 c108 (.A0(net11),
    .A1(net34),
    .A2(net41),
    .A3(net33),
    .S0(net951),
    .S1(net972),
    .X(net44));
 sky130_fd_sc_hd__a2111o_1 c109 (.A1(net41),
    .A2(net38),
    .B1(net44),
    .C1(net7),
    .D1(net43),
    .X(net45));
 sky130_fd_sc_hd__mux4_1 c110 (.A0(net997),
    .A1(net871),
    .A2(net31),
    .A3(net35),
    .S0(net972),
    .S1(net1017),
    .X(net46));
 sky130_fd_sc_hd__and3_1 c111 (.A(net862),
    .B(net6),
    .C(net1006),
    .X(net47));
 sky130_fd_sc_hd__or4bb_1 c112 (.A(net37),
    .B(net6),
    .C_N(net860),
    .D_N(net865),
    .X(net48));
 sky130_fd_sc_hd__and3_2 c113 (.A(net844),
    .B(net862),
    .C(net1020),
    .X(net49));
 sky130_fd_sc_hd__and3_1 c114 (.A(net20),
    .B(net9),
    .C(net37),
    .X(net50));
 sky130_fd_sc_hd__or4bb_2 c115 (.A(net48),
    .B(net46),
    .C_N(net865),
    .D_N(net44),
    .X(net51));
 sky130_fd_sc_hd__or4bb_2 c116 (.A(net990),
    .B(net25),
    .C_N(net50),
    .D_N(net1012),
    .X(net52));
 sky130_fd_sc_hd__and3_1 c117 (.A(net51),
    .B(net48),
    .C(net18),
    .X(net53));
 sky130_fd_sc_hd__and3_2 c118 (.A(net6),
    .B(net50),
    .C(net1017),
    .X(net894));
 sky130_fd_sc_hd__a2111o_1 c119 (.A1(net9),
    .A2(net49),
    .B1(net954),
    .C1(net1045),
    .D1(net1014),
    .X(net54));
 sky130_fd_sc_hd__a2111o_1 c120 (.A1(net1006),
    .A2(net51),
    .B1(net18),
    .C1(net971),
    .D1(net865),
    .X(net55));
 sky130_fd_sc_hd__a2111o_2 c121 (.A1(net18),
    .A2(net25),
    .B1(net55),
    .C1(net51),
    .D1(net954),
    .X(net913));
 sky130_fd_sc_hd__and3_1 c122 (.A(net833),
    .B(net913),
    .C(net49),
    .X(net56));
 sky130_fd_sc_hd__mux4_1 c123 (.A0(net56),
    .A1(net54),
    .A2(net1017),
    .A3(net51),
    .S0(net833),
    .S1(net1045),
    .X(net57));
 sky130_fd_sc_hd__and3_1 c124 (.A(net31),
    .B(net47),
    .C(net954),
    .X(net58));
 sky130_fd_sc_hd__a2111o_1 c125 (.A1(net1014),
    .A2(net55),
    .B1(net47),
    .C1(net954),
    .D1(net58),
    .X(net59));
 sky130_fd_sc_hd__mux4_2 c126 (.A0(net55),
    .A1(net52),
    .A2(net954),
    .A3(net6),
    .S0(net1020),
    .S1(net751),
    .X(net60));
 sky130_fd_sc_hd__mux4_1 c127 (.A0(net871),
    .A1(net51),
    .A2(net60),
    .A3(net9),
    .S0(net1005),
    .S1(net954),
    .X(net61));
 sky130_fd_sc_hd__a2111o_1 c128 (.A1(net60),
    .A2(net48),
    .B1(net954),
    .C1(net59),
    .D1(net973),
    .X(net62));
 sky130_fd_sc_hd__mux4_1 c129 (.A0(net44),
    .A1(net60),
    .A2(net62),
    .A3(net973),
    .S0(net49),
    .S1(net61),
    .X(net63));
 sky130_fd_sc_hd__mux4_1 c130 (.A0(net46),
    .A1(net62),
    .A2(net56),
    .A3(net50),
    .S0(net6),
    .S1(net927),
    .X(net64));
 sky130_fd_sc_hd__sdfbbn_1 c131 (.CLK_N(clknet_4_14_0_clk),
    .D(net60),
    .RESET_B(net61),
    .SCD(net46),
    .SCE(net9),
    .SET_B(net927),
    .Q(net66),
    .Q_N(net65));
 sky130_fd_sc_hd__and3_1 c132 (.A(net1018),
    .B(net1015),
    .C(net995),
    .X(net67));
 sky130_fd_sc_hd__or4bb_4 c133 (.A(net67),
    .B(net703),
    .C_N(net1001),
    .D_N(net1021),
    .X(net68));
 sky130_fd_sc_hd__and3_1 c134 (.A(net1017),
    .B(net996),
    .C(net1021),
    .X(net69));
 sky130_fd_sc_hd__and3_1 c135 (.A(net1001),
    .B(net1004),
    .C(net995),
    .X(net70));
 sky130_fd_sc_hd__and3_2 c136 (.A(net1001),
    .B(net1015),
    .C(net998),
    .X(net71));
 sky130_fd_sc_hd__and3_2 c137 (.A(net995),
    .B(net996),
    .C(net991),
    .X(net72));
 sky130_fd_sc_hd__and3_2 c138 (.A(net1013),
    .B(net1020),
    .C(net67),
    .X(net73));
 sky130_fd_sc_hd__and3_4 c139 (.A(net67),
    .B(net995),
    .C(net991),
    .X(net74));
 sky130_fd_sc_hd__and3_2 c140 (.A(net1024),
    .B(net703),
    .C(net984),
    .X(net75));
 sky130_fd_sc_hd__a2111o_4 c141 (.A1(net983),
    .A2(net995),
    .B1(net1015),
    .C1(net75),
    .D1(net998),
    .X(net76));
 sky130_fd_sc_hd__a2111o_1 c142 (.A1(net1021),
    .A2(net1023),
    .B1(net1001),
    .C1(net983),
    .D1(net991),
    .X(net77));
 sky130_fd_sc_hd__and2_2 c143 (.A(net1011),
    .B(net1024),
    .X(net78));
 sky130_fd_sc_hd__and3_4 c144 (.A(net76),
    .B(net1008),
    .C(net78),
    .X(net79));
 sky130_fd_sc_hd__and3_2 c145 (.A(net993),
    .B(net67),
    .C(net1003),
    .X(net80));
 sky130_fd_sc_hd__and3_4 c146 (.A(net80),
    .B(net1023),
    .C(net980),
    .X(net81));
 sky130_fd_sc_hd__mux4_2 c147 (.A0(net991),
    .A1(net1001),
    .A2(net79),
    .A3(net81),
    .S0(net998),
    .S1(net983),
    .X(net82));
 sky130_fd_sc_hd__and3_1 c148 (.A(net993),
    .B(net969),
    .C(net980),
    .X(net83));
 sky130_fd_sc_hd__mux4_2 c149 (.A0(net80),
    .A1(net1023),
    .A2(net827),
    .A3(net1002),
    .S0(net1004),
    .S1(net71),
    .X(net84));
 sky130_fd_sc_hd__mux4_2 c150 (.A0(net71),
    .A1(net1011),
    .A2(net84),
    .A3(net1008),
    .S0(net980),
    .S1(net74),
    .X(net85));
 sky130_fd_sc_hd__and3_2 c151 (.A(net84),
    .B(net85),
    .C(net67),
    .X(net86));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net85),
    .A1(net83),
    .A2(net983),
    .A3(net84),
    .S0(net79),
    .S1(net86),
    .X(net87));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net87),
    .A1(net84),
    .A2(net85),
    .A3(net86),
    .S0(net994),
    .S1(net1023),
    .X(net88));
 sky130_fd_sc_hd__a2111o_1 c154 (.A1(net847),
    .A2(net78),
    .B1(net1004),
    .C1(net1012),
    .D1(net995),
    .X(net903));
 sky130_fd_sc_hd__and3_2 c155 (.A(net998),
    .B(net86),
    .C(net68),
    .X(net89));
 sky130_fd_sc_hd__and3_1 c156 (.A(net854),
    .B(net1014),
    .C(net84),
    .X(net90));
 sky130_fd_sc_hd__or4bb_4 c157 (.A(net1018),
    .B(net83),
    .C_N(net1012),
    .D_N(net853),
    .X(net91));
 sky130_fd_sc_hd__or4bb_2 c158 (.A(net834),
    .B(net838),
    .C_N(net1009),
    .D_N(net981),
    .X(net92));
 sky130_fd_sc_hd__a2111o_1 c159 (.A1(net90),
    .A2(net836),
    .B1(net827),
    .C1(net969),
    .D1(net1015),
    .X(net93));
 sky130_fd_sc_hd__and3_1 c160 (.A(net838),
    .B(net91),
    .C(net93),
    .X(net94));
 sky130_fd_sc_hd__and3_2 c161 (.A(net93),
    .B(net836),
    .C(net81),
    .X(net95));
 sky130_fd_sc_hd__mux4_2 c162 (.A0(net95),
    .A1(net92),
    .A2(net1013),
    .A3(net837),
    .S0(net981),
    .S1(net998),
    .X(net96));
 sky130_fd_sc_hd__a2111o_2 c163 (.A1(net89),
    .A2(net983),
    .B1(net91),
    .C1(net838),
    .D1(net981),
    .X(net881));
 sky130_fd_sc_hd__a2111o_4 c164 (.A1(net703),
    .A2(net853),
    .B1(net1009),
    .C1(net1002),
    .D1(net95),
    .X(net97));
 sky130_fd_sc_hd__a2111o_4 c165 (.A1(net97),
    .A2(net969),
    .B1(net836),
    .C1(net844),
    .D1(net981),
    .X(net98));
 sky130_fd_sc_hd__a2111o_2 c166 (.A1(net96),
    .A2(net1024),
    .B1(net98),
    .C1(net837),
    .D1(net833),
    .X(net99));
 sky130_fd_sc_hd__a2111o_4 c167 (.A1(net99),
    .A2(net94),
    .B1(net84),
    .C1(net96),
    .D1(net98),
    .X(net100));
 sky130_fd_sc_hd__a2111o_4 c168 (.A1(net89),
    .A2(net100),
    .B1(net92),
    .C1(net1017),
    .D1(net960),
    .X(net101));
 sky130_fd_sc_hd__mux4_2 c169 (.A0(net96),
    .A1(net99),
    .A2(net91),
    .A3(net100),
    .S0(net97),
    .S1(net847),
    .X(net102));
 sky130_fd_sc_hd__a2111o_4 c170 (.A1(net94),
    .A2(net89),
    .B1(net100),
    .C1(net1018),
    .D1(net97),
    .X(net103));
 sky130_fd_sc_hd__a2111o_4 c171 (.A1(net846),
    .A2(net90),
    .B1(net960),
    .C1(net949),
    .D1(net1003),
    .X(net104));
 sky130_fd_sc_hd__mux4_2 c172 (.A0(net102),
    .A1(net100),
    .A2(net827),
    .A3(net104),
    .S0(net97),
    .S1(net949),
    .X(net919));
 sky130_fd_sc_hd__mux4_2 c173 (.A0(net104),
    .A1(net95),
    .A2(net943),
    .A3(net847),
    .S0(net949),
    .S1(net100),
    .X(net105));
 sky130_fd_sc_hd__mux4_2 c174 (.A0(net100),
    .A1(net980),
    .A2(net949),
    .A3(net991),
    .S0(net84),
    .S1(net936),
    .X(net106));
 sky130_fd_sc_hd__mux4_2 c175 (.A0(net936),
    .A1(net841),
    .A2(net106),
    .A3(net943),
    .S0(net961),
    .S1(net104),
    .X(net107));
 sky130_fd_sc_hd__a2111o_1 c176 (.A1(net827),
    .A2(net104),
    .B1(net856),
    .C1(net990),
    .D1(net1022),
    .X(net108));
 sky130_fd_sc_hd__and3_1 c177 (.A(net94),
    .B(net1),
    .C(net1003),
    .X(net914));
 sky130_fd_sc_hd__and3_2 c178 (.A(net83),
    .B(net870),
    .C(net86),
    .X(net109));
 sky130_fd_sc_hd__a2111o_4 c179 (.A1(net869),
    .A2(net106),
    .B1(net991),
    .C1(net847),
    .D1(net998),
    .X(net110));
 sky130_fd_sc_hd__and3_2 c180 (.A(net952),
    .B(net2),
    .C(net1009),
    .X(net111));
 sky130_fd_sc_hd__a2111o_4 c181 (.A1(net1002),
    .A2(net840),
    .B1(net856),
    .C1(net873),
    .D1(net943),
    .X(net112));
 sky130_fd_sc_hd__and3_4 c182 (.A(net844),
    .B(net1),
    .C(net1011),
    .X(net113));
 sky130_fd_sc_hd__and3_1 c183 (.A(net97),
    .B(net858),
    .C(net109),
    .X(net114));
 sky130_fd_sc_hd__a2111o_1 c184 (.A1(net114),
    .A2(net81),
    .B1(net110),
    .C1(net852),
    .D1(net847),
    .X(net115));
 sky130_fd_sc_hd__or4bb_4 c185 (.A(net113),
    .B(net846),
    .C_N(net1001),
    .D_N(net114),
    .X(net116));
 sky130_fd_sc_hd__and3_1 c186 (.A(net79),
    .B(net107),
    .C(net114),
    .X(net117));
 sky130_fd_sc_hd__a2111o_1 c187 (.A1(net849),
    .A2(net870),
    .B1(net113),
    .C1(net116),
    .D1(net995),
    .X(net118));
 sky130_fd_sc_hd__and3_1 c188 (.A(net112),
    .B(net949),
    .C(net991),
    .X(net119));
 sky130_fd_sc_hd__and3_2 c189 (.A(net84),
    .B(net2),
    .C(net952),
    .X(net120));
 sky130_fd_sc_hd__and3_2 c190 (.A(net120),
    .B(net114),
    .C(net119),
    .X(net121));
 sky130_fd_sc_hd__a2111o_1 c191 (.A1(net119),
    .A2(net120),
    .B1(net865),
    .C1(net1009),
    .D1(net1006),
    .X(net122));
 sky130_fd_sc_hd__a2111o_4 c192 (.A1(net116),
    .A2(net114),
    .B1(net935),
    .C1(net1014),
    .D1(net952),
    .X(net123));
 sky130_fd_sc_hd__a2111o_1 c193 (.A1(net935),
    .A2(net117),
    .B1(net119),
    .C1(net121),
    .D1(net108),
    .X(net124));
 sky130_fd_sc_hd__a2111o_4 c194 (.A1(net118),
    .A2(net115),
    .B1(net120),
    .C1(net124),
    .D1(net1007),
    .X(net909));
 sky130_fd_sc_hd__and3_2 c195 (.A(net111),
    .B(net121),
    .C(net935),
    .X(net125));
 sky130_fd_sc_hd__mux4_2 c196 (.A0(net124),
    .A1(net119),
    .A2(net123),
    .A3(net863),
    .S0(net120),
    .S1(net125),
    .X(net126));
 sky130_fd_sc_hd__mux4_2 c197 (.A0(net93),
    .A1(net108),
    .A2(net97),
    .A3(net111),
    .S0(net113),
    .S1(net116),
    .X(net127));
 sky130_fd_sc_hd__and3_1 c198 (.A(net111),
    .B(net74),
    .C(net109),
    .X(net128));
 sky130_fd_sc_hd__and3_4 c199 (.A(net21),
    .B(net79),
    .C(net109),
    .X(net891));
 sky130_fd_sc_hd__and3_4 c200 (.A(net874),
    .B(net868),
    .C(net1007),
    .X(net129));
 sky130_fd_sc_hd__and3_1 c201 (.A(net5),
    .B(net129),
    .C(net992),
    .X(net130));
 sky130_fd_sc_hd__a2111o_1 c202 (.A1(net949),
    .A2(net128),
    .B1(net14),
    .C1(net104),
    .D1(net1029),
    .X(net131));
 sky130_fd_sc_hd__a2111o_2 c203 (.A1(net106),
    .A2(net124),
    .B1(net1038),
    .C1(net130),
    .D1(net849),
    .X(net132));
 sky130_fd_sc_hd__a2111o_1 c204 (.A1(net103),
    .A2(net833),
    .B1(net129),
    .C1(net1044),
    .D1(net1000),
    .X(net133));
 sky130_fd_sc_hd__and3_2 c205 (.A(net845),
    .B(net115),
    .C(net0),
    .X(net134));
 sky130_fd_sc_hd__a2111o_1 c206 (.A1(net74),
    .A2(net134),
    .B1(net842),
    .C1(net1044),
    .D1(net81),
    .X(net135));
 sky130_fd_sc_hd__mux4_1 c207 (.A0(net14),
    .A1(net113),
    .A2(net134),
    .A3(net103),
    .S0(net991),
    .S1(net1038),
    .X(net136));
 sky130_fd_sc_hd__and3_1 c208 (.A(net130),
    .B(net79),
    .C(net20),
    .X(net137));
 sky130_fd_sc_hd__and3_1 c209 (.A(net129),
    .B(net863),
    .C(net957),
    .X(net138));
 sky130_fd_sc_hd__sdfbbn_2 c210 (.CLK_N(clknet_4_10_0_clk),
    .D(net134),
    .RESET_B(net874),
    .SCD(net957),
    .SCE(net136),
    .SET_B(net132),
    .Q(net888),
    .Q_N(net139));
 sky130_fd_sc_hd__mux4_2 c211 (.A0(net842),
    .A1(net112),
    .A2(net123),
    .A3(net1009),
    .S0(net971),
    .S1(net957),
    .X(net140));
 sky130_fd_sc_hd__a2111o_1 c212 (.A1(net841),
    .A2(net138),
    .B1(net140),
    .C1(net958),
    .D1(net952),
    .X(net141));
 sky130_fd_sc_hd__mux4_2 c213 (.A0(net133),
    .A1(net20),
    .A2(net5),
    .A3(net14),
    .S0(net24),
    .S1(net140),
    .X(net142));
 sky130_fd_sc_hd__mux4_1 c214 (.A0(net128),
    .A1(net132),
    .A2(net1079),
    .A3(net14),
    .S0(net123),
    .S1(net957),
    .X(net143));
 sky130_fd_sc_hd__mux4_1 c215 (.A0(net141),
    .A1(net1033),
    .A2(net142),
    .A3(net957),
    .S0(net983),
    .S1(net111),
    .X(net144));
 sky130_fd_sc_hd__a2111o_1 c216 (.A1(net140),
    .A2(net837),
    .B1(net957),
    .C1(net1044),
    .D1(net753),
    .X(net145));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(net135),
    .A1(net957),
    .A2(net142),
    .A3(net133),
    .S0(net1079),
    .S1(net1049),
    .X(net146));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(net145),
    .A1(net1079),
    .A2(net891),
    .A3(net23),
    .S0(net957),
    .S1(net753),
    .X(net147));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net136),
    .A1(net10),
    .A2(net142),
    .A3(net1009),
    .S0(net111),
    .S1(net989),
    .X(net148));
 sky130_fd_sc_hd__a2111o_4 c220 (.A1(net972),
    .A2(net140),
    .B1(net26),
    .C1(net138),
    .D1(net981),
    .X(net880));
 sky130_fd_sc_hd__sdfbbp_1 c221 (.CLK(clknet_4_11_0_clk),
    .D(net141),
    .RESET_B(net1007),
    .SCD(net37),
    .SCE(net1041),
    .SET_B(net32),
    .Q(net898),
    .Q_N(net149));
 sky130_fd_sc_hd__a2111o_2 c222 (.A1(net958),
    .A2(net943),
    .B1(net972),
    .C1(net989),
    .D1(net754),
    .X(net150));
 sky130_fd_sc_hd__sdfbbn_1 c223 (.CLK_N(clknet_4_14_0_clk),
    .D(net45),
    .RESET_B(net142),
    .SCD(net109),
    .SCE(net1000),
    .SET_B(net68),
    .Q(net152),
    .Q_N(net151));
 sky130_fd_sc_hd__mux4_1 c224 (.A0(net124),
    .A1(net1082),
    .A2(net109),
    .A3(net149),
    .S0(net831),
    .S1(net753),
    .X(net153));
 sky130_fd_sc_hd__a2111o_4 c225 (.A1(net951),
    .A2(net884),
    .B1(net664),
    .C1(net754),
    .D1(net755),
    .X(net154));
 sky130_fd_sc_hd__mux4_2 c226 (.A0(net32),
    .A1(net150),
    .A2(net898),
    .A3(net154),
    .S0(net2),
    .S1(net755),
    .X(net155));
 sky130_fd_sc_hd__mux4_1 c227 (.A0(net27),
    .A1(net874),
    .A2(net1014),
    .A3(net997),
    .S0(net664),
    .S1(net755),
    .X(net156));
 sky130_fd_sc_hd__mux4_1 c228 (.A0(net24),
    .A1(net26),
    .A2(net101),
    .A3(net943),
    .S0(net1000),
    .S1(net755),
    .X(net157));
 sky130_fd_sc_hd__mux4_1 c229 (.A0(net43),
    .A1(net150),
    .A2(net16),
    .A3(net101),
    .S0(net1012),
    .S1(net972),
    .X(net158));
 sky130_fd_sc_hd__a2111o_1 c230 (.A1(net117),
    .A2(net129),
    .B1(net1035),
    .C1(net45),
    .D1(net151),
    .X(net159));
 sky130_fd_sc_hd__mux4_1 c231 (.A0(net113),
    .A1(net960),
    .A2(net863),
    .A3(net149),
    .S0(net1023),
    .S1(net957),
    .X(net160));
 sky130_fd_sc_hd__a2111o_1 c232 (.A1(net156),
    .A2(net40),
    .B1(net26),
    .C1(net1007),
    .D1(net754),
    .X(net161));
 sky130_fd_sc_hd__sdfbbn_2 c233 (.CLK_N(clknet_4_15_0_clk),
    .D(net161),
    .RESET_B(net142),
    .SCD(net116),
    .SCE(net981),
    .SET_B(net754),
    .Q(net904),
    .Q_N(net162));
 sky130_fd_sc_hd__a2111o_1 c234 (.A1(net157),
    .A2(net42),
    .B1(net943),
    .C1(net834),
    .D1(net1081),
    .X(net163));
 sky130_fd_sc_hd__mux4_1 c235 (.A0(net158),
    .A1(net140),
    .A2(net162),
    .A3(net151),
    .S0(net113),
    .S1(net154),
    .X(net164));
 sky130_fd_sc_hd__mux4_2 c236 (.A0(net155),
    .A1(net149),
    .A2(net162),
    .A3(net156),
    .S0(net664),
    .X(net674));
 sky130_fd_sc_hd__mux4_1 c237 (.A0(net2),
    .A1(net150),
    .A2(net904),
    .A3(net27),
    .S0(net837),
    .S1(net113),
    .X(net166));
 sky130_fd_sc_hd__mux4_1 c238 (.A0(net166),
    .A1(net838),
    .A2(net158),
    .A3(net164),
    .S0(net1010),
    .S1(net162),
    .X(net167));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net164),
    .A1(net113),
    .A2(net166),
    .A3(net24),
    .S0(net35),
    .S1(net675),
    .X(net168));
 sky130_fd_sc_hd__mux4_1 c240 (.A0(net1035),
    .A1(net904),
    .A2(net161),
    .A3(net1083),
    .S0(net117),
    .S1(net675),
    .X(net169));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(net115),
    .A1(net26),
    .A2(net868),
    .A3(net15),
    .S0(net756),
    .S1(clknet_1_1__leaf_net758),
    .X(net170));
 sky130_fd_sc_hd__mux4_2 c242 (.A0(net834),
    .A1(net50),
    .A2(net25),
    .A3(net1014),
    .S0(net674),
    .S1(net751),
    .X(net171));
 sky130_fd_sc_hd__mux4_2 c243 (.A0(net865),
    .A1(net54),
    .A2(net898),
    .A3(net1023),
    .S0(net971),
    .S1(net25),
    .X(net885));
 sky130_fd_sc_hd__mux4_1 c244 (.A0(net854),
    .A1(net160),
    .A2(net139),
    .A3(net31),
    .S0(net931),
    .S1(net1041),
    .X(net172));
 sky130_fd_sc_hd__sdfbbp_1 c245 (.CLK(clknet_4_11_0_clk),
    .D(net913),
    .RESET_B(net931),
    .SCD(net29),
    .SCE(net674),
    .SET_B(clknet_1_0__leaf_net759),
    .Q(net174),
    .Q_N(net173));
 sky130_fd_sc_hd__mux4_1 c246 (.A0(net860),
    .A1(net981),
    .A2(net149),
    .A3(net909),
    .S0(net138),
    .S1(clknet_1_0__leaf_net759),
    .X(net175));
 sky130_fd_sc_hd__mux4_1 c247 (.A0(net61),
    .A1(net1037),
    .A2(net1020),
    .A3(net880),
    .S1(clknet_1_1__leaf_net759),
    .X(net709));
 sky130_fd_sc_hd__mux4_1 c248 (.A0(net138),
    .A1(net943),
    .A2(net173),
    .A3(net992),
    .S0(net1022),
    .S1(clknet_1_0__leaf_net759),
    .X(net905));
 sky130_fd_sc_hd__mux4_1 c249 (.A0(net174),
    .A1(net53),
    .A2(net49),
    .A3(net25),
    .S0(net1017),
    .S1(clknet_1_0__leaf_net759),
    .X(net924));
 sky130_fd_sc_hd__mux4_2 c250 (.A0(net29),
    .A1(clknet_1_0__leaf_net905),
    .A2(net1037),
    .A3(net52),
    .S0(net898),
    .S1(net112),
    .X(net902));
 sky130_fd_sc_hd__mux4_2 c251 (.A0(net25),
    .A1(net157),
    .A2(net59),
    .A3(clknet_1_0__leaf_net902),
    .S0(clknet_1_1__leaf_net905),
    .S1(clknet_1_0__leaf_net709),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 c252 (.A0(net833),
    .A1(clknet_1_0__leaf_net905),
    .A2(net20),
    .A3(net1080),
    .S0(net954),
    .S1(net981),
    .X(net178));
 sky130_fd_sc_hd__mux4_1 c253 (.A0(net54),
    .A1(net885),
    .A2(net20),
    .A3(net1045),
    .S0(net981),
    .S1(clknet_1_0__leaf_net901),
    .X(net179));
 sky130_fd_sc_hd__mux4_2 c254 (.A0(clknet_1_1__leaf_net179),
    .A1(net982),
    .A2(net60),
    .A3(net835),
    .S0(clknet_1_1__leaf_net709),
    .S1(clknet_1_1__leaf_net759),
    .X(net180));
 sky130_fd_sc_hd__mux4_1 c255 (.A0(net160),
    .A1(net60),
    .A2(net860),
    .A3(net943),
    .S0(net960),
    .S1(clknet_1_0__leaf_net901),
    .X(net910));
 sky130_fd_sc_hd__mux4_1 c256 (.A0(net47),
    .A1(clknet_1_0__leaf_net177),
    .A2(clknet_1_0__leaf_net924),
    .A3(clknet_1_0__leaf_net180),
    .S0(clknet_1_0__leaf_net910),
    .S1(clknet_1_0__leaf_net901),
    .X(net181));
 sky130_fd_sc_hd__mux4_1 c257 (.A0(net35),
    .A1(net62),
    .A2(net1040),
    .A3(net60),
    .S0(net1023),
    .S1(clknet_1_1__leaf_net901),
    .X(net182));
 sky130_fd_sc_hd__mux4_2 c258 (.A0(net59),
    .A1(clknet_1_0__leaf_net180),
    .A2(net884),
    .A3(net952),
    .S0(net52),
    .S1(clknet_1_1__leaf_net901),
    .X(net183));
 sky130_fd_sc_hd__mux4_1 c259 (.A0(clknet_1_1__leaf_net177),
    .A1(net973),
    .A2(net29),
    .A3(net702),
    .S0(net899),
    .S1(clknet_1_1__leaf_net759),
    .X(net184));
 sky130_fd_sc_hd__mux4_2 c260 (.A0(net171),
    .A1(net58),
    .A2(net65),
    .A3(net173),
    .S0(net749),
    .S1(clknet_1_0__leaf_net759),
    .X(net185));
 sky130_fd_sc_hd__mux4_2 c261 (.A0(net1017),
    .A1(net185),
    .A2(net952),
    .A3(net749),
    .S0(clknet_1_0__leaf_net759),
    .S1(clknet_1_0__leaf_net901),
    .X(net186));
 sky130_fd_sc_hd__mux4_2 c262 (.A0(clknet_1_0__leaf_net186),
    .A1(net112),
    .A2(net854),
    .A3(net174),
    .S0(net749),
    .S1(clknet_1_0__leaf_net901),
    .X(net187));
 sky130_fd_sc_hd__mux4_2 c263 (.A0(clknet_1_0__leaf_net177),
    .A1(net187),
    .A2(clknet_1_1__leaf_net186),
    .A3(clknet_1_1__leaf_net905),
    .S0(net885),
    .S1(clknet_1_0__leaf_net759),
    .X(net188));
 sky130_fd_sc_hd__and3_1 c264 (.A(net1023),
    .B(net993),
    .C(net980),
    .X(net189));
 sky130_fd_sc_hd__and3_2 c265 (.A(net1015),
    .B(net1002),
    .C(net978),
    .X(net190));
 sky130_fd_sc_hd__and3_4 c266 (.A(net998),
    .B(net976),
    .C(net1015),
    .X(net191));
 sky130_fd_sc_hd__and3_4 c267 (.A(net976),
    .B(net74),
    .C(net998),
    .X(net192));
 sky130_fd_sc_hd__a2111o_4 c268 (.A1(net81),
    .A2(net74),
    .B1(net191),
    .C1(net1008),
    .D1(net977),
    .X(net193));
 sky130_fd_sc_hd__and3_2 c269 (.A(net77),
    .B(net87),
    .C(net976),
    .X(net194));
 sky130_fd_sc_hd__a2111o_2 c270 (.A1(net1024),
    .A2(net75),
    .B1(net703),
    .C1(net977),
    .D1(net1004),
    .X(net195));
 sky130_fd_sc_hd__and3_2 c271 (.A(net193),
    .B(net703),
    .C(net977),
    .X(net196));
 sky130_fd_sc_hd__and3_4 c272 (.A(net827),
    .B(net974),
    .C(net976),
    .X(net197));
 sky130_fd_sc_hd__and3_2 c273 (.A(net67),
    .B(net191),
    .C(net977),
    .X(net198));
 sky130_fd_sc_hd__and3_2 c274 (.A(net193),
    .B(net192),
    .C(net984),
    .X(net199));
 sky130_fd_sc_hd__a2111o_4 c275 (.A1(net974),
    .A2(net78),
    .B1(net191),
    .C1(net967),
    .D1(net976),
    .X(net200));
 sky130_fd_sc_hd__or4bb_1 c276 (.A(net196),
    .B(net961),
    .C_N(net68),
    .D_N(net976),
    .X(net201));
 sky130_fd_sc_hd__and3_2 c277 (.A(net1024),
    .B(net974),
    .C(net1013),
    .X(net202));
 sky130_fd_sc_hd__and3_1 c278 (.A(net202),
    .B(net198),
    .C(net197),
    .X(net203));
 sky130_fd_sc_hd__and3_1 c279 (.A(net201),
    .B(net78),
    .C(net963),
    .X(net204));
 sky130_fd_sc_hd__mux4_2 c280 (.A0(net192),
    .A1(net995),
    .A2(net974),
    .A3(net976),
    .S0(net196),
    .S1(net197),
    .X(net205));
 sky130_fd_sc_hd__mux4_2 c281 (.A0(net204),
    .A1(net202),
    .A2(net78),
    .A3(net967),
    .S0(net974),
    .S1(net963),
    .X(net206));
 sky130_fd_sc_hd__mux4_2 c282 (.A0(net1003),
    .A1(net197),
    .A2(net202),
    .A3(net963),
    .S0(net998),
    .S1(net976),
    .X(net207));
 sky130_fd_sc_hd__mux4_2 c283 (.A0(net194),
    .A1(net201),
    .A2(net703),
    .A3(net198),
    .S0(net963),
    .S1(net976),
    .X(net208));
 sky130_fd_sc_hd__mux4_2 c284 (.A0(net974),
    .A1(net205),
    .A2(net198),
    .A3(net204),
    .S0(net964),
    .S1(net976),
    .X(net209));
 sky130_fd_sc_hd__mux4_2 c285 (.A0(net208),
    .A1(net205),
    .A2(net209),
    .A3(net192),
    .S0(net974),
    .S1(net1003),
    .X(net210));
 sky130_fd_sc_hd__and3_1 c286 (.A(net107),
    .B(net840),
    .C(net207),
    .X(net906));
 sky130_fd_sc_hd__or4bb_4 c287 (.A(net1022),
    .B(net198),
    .C_N(net1003),
    .D_N(net853),
    .X(net211));
 sky130_fd_sc_hd__or4bb_2 c288 (.A(net1009),
    .B(net208),
    .C_N(net949),
    .D_N(net206),
    .X(net917));
 sky130_fd_sc_hd__or4bb_4 c289 (.A(net194),
    .B(net103),
    .C_N(net962),
    .D_N(net964),
    .X(net212));
 sky130_fd_sc_hd__a2111o_4 c290 (.A1(net92),
    .A2(net87),
    .B1(net91),
    .C1(net1009),
    .D1(net977),
    .X(net213));
 sky130_fd_sc_hd__a2111o_2 c291 (.A1(net90),
    .A2(net827),
    .B1(net967),
    .C1(net961),
    .D1(net106),
    .X(net214));
 sky130_fd_sc_hd__and3_1 c292 (.A(net106),
    .B(net944),
    .C(net943),
    .X(net215));
 sky130_fd_sc_hd__or4bb_2 c293 (.A(net215),
    .B(net214),
    .C_N(net995),
    .D_N(net933),
    .X(net216));
 sky130_fd_sc_hd__and3_4 c294 (.A(net962),
    .B(net104),
    .C(net974),
    .X(net217));
 sky130_fd_sc_hd__a2111o_2 c295 (.A1(net83),
    .A2(net1009),
    .B1(net991),
    .C1(net964),
    .D1(net213),
    .X(net218));
 sky130_fd_sc_hd__or4bb_4 c296 (.A(net944),
    .B(net214),
    .C_N(net213),
    .D_N(net217),
    .X(net219));
 sky130_fd_sc_hd__or4bb_1 c297 (.A(net78),
    .B(net853),
    .C_N(net962),
    .D_N(net208),
    .X(net220));
 sky130_fd_sc_hd__a2111o_1 c298 (.A1(net213),
    .A2(net71),
    .B1(net96),
    .C1(net216),
    .D1(net944),
    .X(net221));
 sky130_fd_sc_hd__or4bb_4 c299 (.A(net832),
    .B(net217),
    .C_N(net219),
    .D_N(net1024),
    .X(net222));
 sky130_fd_sc_hd__or4bb_2 c300 (.A(net222),
    .B(net214),
    .C_N(net936),
    .D_N(net948),
    .X(net223));
 sky130_fd_sc_hd__and3_1 c301 (.A(net222),
    .B(net102),
    .C(net950),
    .X(net224));
 sky130_fd_sc_hd__or4bb_2 c302 (.A(net86),
    .B(net218),
    .C_N(net219),
    .D_N(net950),
    .X(net225));
 sky130_fd_sc_hd__a2111o_1 c303 (.A1(net219),
    .A2(net224),
    .B1(net834),
    .C1(net950),
    .D1(net192),
    .X(net226));
 sky130_fd_sc_hd__mux4_2 c304 (.A0(net225),
    .A1(net213),
    .A2(net222),
    .A3(net1012),
    .S0(net96),
    .S1(net102),
    .X(net227));
 sky130_fd_sc_hd__mux4_1 c305 (.A0(net227),
    .A1(net832),
    .A2(net222),
    .A3(net950),
    .S0(net202),
    .S1(net962),
    .X(net228));
 sky130_fd_sc_hd__mux4_1 c306 (.A0(net102),
    .A1(net223),
    .A2(net933),
    .A3(net213),
    .S0(net962),
    .S1(net227),
    .X(net229));
 sky130_fd_sc_hd__mux4_1 c307 (.A0(net86),
    .A1(net227),
    .A2(net933),
    .A3(net202),
    .S0(net676),
    .S1(net988),
    .X(net230));
 sky130_fd_sc_hd__mux4_2 c308 (.A0(net71),
    .A1(net108),
    .A2(net193),
    .A3(net106),
    .S0(net984),
    .S1(net219),
    .X(net231));
 sky130_fd_sc_hd__or4bb_1 c309 (.A(net840),
    .B(net104),
    .C_N(net849),
    .D_N(net1006),
    .X(net892));
 sky130_fd_sc_hd__a2111o_4 c310 (.A1(net865),
    .A2(net123),
    .B1(net936),
    .C1(net1012),
    .D1(net999),
    .X(net889));
 sky130_fd_sc_hd__mux4_1 c311 (.A0(net78),
    .A1(net120),
    .A2(net917),
    .A3(net119),
    .S0(net106),
    .S1(net941),
    .X(net232));
 sky130_fd_sc_hd__or4bb_2 c312 (.A(net191),
    .B(net889),
    .C_N(net835),
    .D_N(net941),
    .X(net233));
 sky130_fd_sc_hd__or4bb_1 c313 (.A(net233),
    .B(net889),
    .C_N(net960),
    .D_N(net194),
    .X(net234));
 sky130_fd_sc_hd__or4bb_1 c314 (.A(net119),
    .B(net79),
    .C_N(net223),
    .X(net235));
 sky130_fd_sc_hd__or4bb_4 c315 (.A(net967),
    .B(net118),
    .C_N(net110),
    .D_N(net127),
    .X(net236));
 sky130_fd_sc_hd__a2111o_1 c316 (.A1(net108),
    .A2(net233),
    .B1(net218),
    .C1(net941),
    .D1(net745),
    .X(net237));
 sky130_fd_sc_hd__sdfbbn_2 c317 (.CLK_N(clknet_4_8_0_clk),
    .D(net118),
    .RESET_B(net227),
    .SCD(net125),
    .SCE(net889),
    .SET_B(net941),
    .Q(net239),
    .Q_N(net238));
 sky130_fd_sc_hd__a2111o_1 c318 (.A1(net236),
    .A2(net73),
    .B1(net197),
    .C1(net1006),
    .D1(net745),
    .X(net240));
 sky130_fd_sc_hd__a2111o_2 c319 (.A1(net225),
    .A2(net832),
    .B1(net996),
    .C1(net238),
    .D1(net745),
    .X(net241));
 sky130_fd_sc_hd__a2111o_4 c320 (.A1(net91),
    .A2(net71),
    .B1(net840),
    .C1(net193),
    .D1(net110),
    .X(net242));
 sky130_fd_sc_hd__mux4_1 c321 (.A0(net127),
    .A1(net873),
    .A2(net233),
    .A3(net863),
    .S0(net242),
    .S1(net745),
    .X(net243));
 sky130_fd_sc_hd__or4bb_1 c322 (.A(net232),
    .B(net233),
    .C_N(net236),
    .D_N(net209),
    .X(net244));
 sky130_fd_sc_hd__a2111o_1 c323 (.A1(net221),
    .A2(net982),
    .B1(net126),
    .C1(net222),
    .D1(net727),
    .X(net245));
 sky130_fd_sc_hd__or4bb_4 c324 (.A(net847),
    .B(net964),
    .C_N(net684),
    .D_N(net745),
    .X(net246));
 sky130_fd_sc_hd__mux4_2 c325 (.A0(net827),
    .A1(net239),
    .A2(net933),
    .A3(net246),
    .S0(net236),
    .S1(net727),
    .X(net247));
 sky130_fd_sc_hd__a2111o_4 c326 (.A1(net247),
    .A2(net231),
    .B1(net849),
    .C1(net1031),
    .D1(net699),
    .X(net248));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(net120),
    .A1(net248),
    .A2(net214),
    .A3(net238),
    .S0(net889),
    .S1(net236),
    .X(net249));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(net248),
    .A1(net238),
    .A2(net127),
    .A3(net242),
    .S0(net233),
    .S1(net721),
    .X(net250));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net121),
    .A1(net232),
    .A2(net248),
    .A3(net988),
    .S1(net727),
    .X(net251));
 sky130_fd_sc_hd__a2111o_1 c330 (.A1(net1031),
    .A2(net194),
    .B1(net248),
    .C1(net935),
    .D1(net79),
    .X(net252));
 sky130_fd_sc_hd__mux4_1 c331 (.A0(net109),
    .A1(net106),
    .A2(net248),
    .A3(net962),
    .S0(net868),
    .S1(net834),
    .X(net253));
 sky130_fd_sc_hd__a2111o_1 c332 (.A1(net79),
    .A2(net1038),
    .B1(net1044),
    .C1(net842),
    .D1(net974),
    .X(net254));
 sky130_fd_sc_hd__mux4_1 c333 (.A0(net240),
    .A1(net142),
    .A2(net16),
    .A3(net949),
    .S0(net827),
    .S1(net761),
    .X(net255));
 sky130_fd_sc_hd__a2111o_1 c334 (.A1(net223),
    .A2(net129),
    .B1(net240),
    .C1(net122),
    .D1(net760),
    .X(net256));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(net1038),
    .A1(net917),
    .A2(net198),
    .A3(net82),
    .S0(net1022),
    .S1(net664),
    .X(net257));
 sky130_fd_sc_hd__mux4_1 c336 (.A0(net214),
    .A1(net1038),
    .A2(net941),
    .A3(net677),
    .S0(net721),
    .S1(net761),
    .X(net258));
 sky130_fd_sc_hd__mux4_2 c337 (.A0(net104),
    .A1(net991),
    .A2(net198),
    .A3(net857),
    .S0(net721),
    .S1(net761),
    .X(net259));
 sky130_fd_sc_hd__mux4_1 c338 (.A0(net254),
    .A1(net1009),
    .A2(net1),
    .A3(net122),
    .S0(net79),
    .S1(net145),
    .X(net260));
 sky130_fd_sc_hd__mux4_2 c339 (.A0(net257),
    .A1(net19),
    .A2(net1011),
    .A3(net823),
    .S0(net664),
    .S1(net989),
    .X(net261));
 sky130_fd_sc_hd__mux4_2 c340 (.A0(net214),
    .A1(net212),
    .A2(net211),
    .A3(net257),
    .S0(net19),
    .S1(net714),
    .X(net262));
 sky130_fd_sc_hd__a2111o_2 c341 (.A1(net1001),
    .A2(net1027),
    .B1(net867),
    .C1(net10),
    .D1(net899),
    .X(net263));
 sky130_fd_sc_hd__mux4_2 c342 (.A0(net86),
    .A1(net254),
    .A2(net891),
    .A3(net257),
    .S0(net957),
    .S1(net760),
    .X(net264));
 sky130_fd_sc_hd__mux4_1 c343 (.A0(net132),
    .A1(net967),
    .A2(net264),
    .A3(net130),
    .S0(net664),
    .S1(net677),
    .X(net265));
 sky130_fd_sc_hd__mux4_2 c344 (.A0(net123),
    .A1(net262),
    .A2(net830),
    .A3(net261),
    .S0(net989),
    .S1(net732),
    .X(net266));
 sky130_fd_sc_hd__a2111o_4 c345 (.A1(net123),
    .A2(net891),
    .B1(net259),
    .C1(net139),
    .D1(net721),
    .X(net267));
 sky130_fd_sc_hd__mux4_2 c346 (.A0(net123),
    .A1(net259),
    .A2(net207),
    .A3(net677),
    .S0(net745),
    .S1(net760),
    .X(net268));
 sky130_fd_sc_hd__mux4_2 c347 (.A0(net198),
    .A1(net109),
    .A2(net267),
    .A3(net941),
    .S0(net264),
    .S1(net899),
    .X(net269));
 sky130_fd_sc_hd__mux4_2 c348 (.A0(net259),
    .A1(net109),
    .A2(net254),
    .A3(net121),
    .S0(net857),
    .S1(net899),
    .X(net270));
 sky130_fd_sc_hd__mux4_2 c349 (.A0(net130),
    .A1(net1012),
    .A2(net270),
    .A3(net267),
    .S0(net258),
    .S1(net714),
    .X(net271));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(net258),
    .A1(net240),
    .A2(net262),
    .A3(net86),
    .S0(net958),
    .S1(net271),
    .X(net272));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net264),
    .A1(net270),
    .A2(net936),
    .A3(net132),
    .S0(net664),
    .S1(net1065),
    .X(net273));
 sky130_fd_sc_hd__mux4_1 c352 (.A0(net135),
    .A1(net248),
    .A2(net271),
    .A3(net1045),
    .S0(net88),
    .S1(net760),
    .X(net274));
 sky130_fd_sc_hd__mux4_1 c353 (.A0(net39),
    .A1(net823),
    .A2(net42),
    .A3(net129),
    .S0(net212),
    .S1(net731),
    .X(net275));
 sky130_fd_sc_hd__mux4_1 c354 (.A0(clknet_1_0__leaf_net170),
    .A1(net857),
    .A2(net992),
    .A3(net823),
    .S0(net958),
    .S1(clknet_1_0__leaf_net758),
    .X(net276));
 sky130_fd_sc_hd__mux4_1 c355 (.A0(net40),
    .A1(net831),
    .A2(net865),
    .A3(net269),
    .S0(net264),
    .S1(net942),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 c356 (.A0(net152),
    .A1(net246),
    .A2(net264),
    .A3(net972),
    .S0(clknet_1_1__leaf_net170),
    .S1(net734),
    .X(net916));
 sky130_fd_sc_hd__mux4_1 c357 (.A0(net246),
    .A1(net152),
    .A2(net969),
    .A3(net865),
    .S0(net731),
    .S1(net762),
    .X(net278));
 sky130_fd_sc_hd__mux4_1 c358 (.A0(net42),
    .A1(net134),
    .A2(net868),
    .A3(net856),
    .S0(net1005),
    .S1(net1070),
    .X(net279));
 sky130_fd_sc_hd__mux4_2 c359 (.A0(net1039),
    .A1(net134),
    .A2(net993),
    .A3(net1023),
    .S0(net955),
    .S1(net1006),
    .X(net923));
 sky130_fd_sc_hd__mux4_1 c360 (.A0(net966),
    .A1(net211),
    .A2(net866),
    .A3(net891),
    .S0(net955),
    .S1(net944),
    .X(net280));
 sky130_fd_sc_hd__mux4_1 c361 (.A0(net33),
    .A1(net280),
    .A2(net1003),
    .A3(net955),
    .S0(clknet_1_1__leaf_net758),
    .S1(net762),
    .X(net281));
 sky130_fd_sc_hd__mux4_1 c362 (.A0(net858),
    .A1(net275),
    .A2(net193),
    .A3(net279),
    .S0(net956),
    .S1(net1051),
    .X(net282));
 sky130_fd_sc_hd__mux4_1 c363 (.A0(net37),
    .A1(net152),
    .A2(net1010),
    .A3(net955),
    .S0(net271),
    .S1(net930),
    .X(net283));
 sky130_fd_sc_hd__mux4_2 c364 (.A0(net150),
    .A1(net225),
    .A2(net993),
    .A3(net1000),
    .S0(net955),
    .S1(net872),
    .X(net284));
 sky130_fd_sc_hd__mux4_1 c365 (.A0(net193),
    .A1(net1011),
    .A2(net955),
    .A3(net713),
    .S0(clknet_1_1__leaf_net758),
    .S1(net920),
    .X(net285));
 sky130_fd_sc_hd__mux4_1 c366 (.A0(clknet_1_1__leaf_net276),
    .A1(net39),
    .A2(net889),
    .A3(net1010),
    .S0(net919),
    .S1(net721),
    .X(net286));
 sky130_fd_sc_hd__mux4_1 c367 (.A0(net1035),
    .A1(net150),
    .A2(net844),
    .A3(net1039),
    .S0(net692),
    .S1(net713),
    .X(net287));
 sky130_fd_sc_hd__mux4_1 c368 (.A0(net142),
    .A1(net285),
    .A2(net956),
    .A3(net212),
    .S0(net756),
    .S1(net763),
    .X(net288));
 sky130_fd_sc_hd__a2111o_2 c369 (.A1(net121),
    .A2(net956),
    .B1(net275),
    .C1(net692),
    .D1(net764),
    .X(net918));
 sky130_fd_sc_hd__mux4_2 c370 (.A0(net205),
    .A1(net837),
    .A2(net918),
    .A3(net956),
    .S0(net925),
    .S1(net764),
    .X(net912));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(clknet_1_1__leaf_net281),
    .A1(net918),
    .A2(net40),
    .A3(net30),
    .S0(net731),
    .S1(net764),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net1036),
    .A1(net31),
    .A2(net923),
    .A3(net247),
    .S0(net713),
    .S1(net1057),
    .X(net290));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net289),
    .A1(net263),
    .A2(net956),
    .A3(net39),
    .S0(net861),
    .S1(net764),
    .X(net911));
 sky130_fd_sc_hd__mux4_1 c374 (.A0(net145),
    .A1(clknet_1_0__leaf_net902),
    .A2(net271),
    .A3(net834),
    .S0(net134),
    .S1(net702),
    .X(net291));
 sky130_fd_sc_hd__mux4_1 c375 (.A0(net66),
    .A1(net856),
    .A2(net861),
    .A3(clknet_1_0__leaf_net179),
    .S0(net974),
    .S1(net952),
    .X(net292));
 sky130_fd_sc_hd__mux4_1 c376 (.A0(net49),
    .A1(net134),
    .A2(net36),
    .A3(net888),
    .S0(net997),
    .S1(net835),
    .X(net293));
 sky130_fd_sc_hd__mux4_1 c377 (.A0(net50),
    .A1(net880),
    .A2(net162),
    .A3(clknet_1_1__leaf_net177),
    .S0(net848),
    .S1(net702),
    .X(net294));
 sky130_fd_sc_hd__mux4_1 c378 (.A0(net271),
    .A1(clknet_1_1__leaf_net180),
    .A2(net960),
    .A3(net898),
    .S0(net997),
    .S1(net925),
    .X(net295));
 sky130_fd_sc_hd__mux4_1 c379 (.A0(net262),
    .A1(net56),
    .A2(net975),
    .A3(net992),
    .S0(net752),
    .S1(clknet_1_0__leaf_net901),
    .X(net296));
 sky130_fd_sc_hd__mux4_1 c380 (.A0(net264),
    .A1(net982),
    .A2(net992),
    .A3(net844),
    .S0(net972),
    .S1(net927),
    .X(net297));
 sky130_fd_sc_hd__mux4_1 c381 (.A0(net868),
    .A1(net297),
    .A2(net271),
    .A3(net952),
    .S0(net899),
    .S1(net748),
    .X(net298));
 sky130_fd_sc_hd__mux4_1 c382 (.A0(net53),
    .A1(net31),
    .A2(net889),
    .A3(net65),
    .S0(clknet_1_1__leaf_net759),
    .S1(net765),
    .X(net299));
 sky130_fd_sc_hd__mux4_1 c383 (.A0(net1023),
    .A1(net270),
    .A2(net884),
    .A3(net1007),
    .S0(net65),
    .S1(net992),
    .X(net300));
 sky130_fd_sc_hd__mux4_1 c384 (.A0(net300),
    .A1(net913),
    .A2(net1040),
    .A3(net284),
    .S0(clknet_1_0__leaf_net709),
    .S1(net748),
    .X(net301));
 sky130_fd_sc_hd__mux4_1 c385 (.A0(clknet_1_0__leaf_net179),
    .A1(net973),
    .A2(net904),
    .A3(net954),
    .S0(net752),
    .S1(net766),
    .X(net302));
 sky130_fd_sc_hd__mux4_1 c386 (.A0(net302),
    .A1(net31),
    .A2(net1020),
    .A3(net1081),
    .S0(net988),
    .S1(net763),
    .X(net303));
 sky130_fd_sc_hd__mux4_1 c387 (.A0(net36),
    .A1(net264),
    .A2(net953),
    .A3(net975),
    .S0(net897),
    .S1(net765),
    .X(net304));
 sky130_fd_sc_hd__mux4_1 c388 (.A0(net299),
    .A1(net953),
    .A2(net37),
    .A3(net877),
    .S0(net749),
    .S1(net766),
    .X(net305));
 sky130_fd_sc_hd__mux4_1 c389 (.A0(net975),
    .A1(net825),
    .A2(net139),
    .A3(net748),
    .S0(net752),
    .S1(clknet_1_1__leaf_net759),
    .X(net306));
 sky130_fd_sc_hd__mux4_1 c390 (.A0(net52),
    .A1(net973),
    .A2(net953),
    .A3(net702),
    .S0(net762),
    .S1(net765),
    .X(net307));
 sky130_fd_sc_hd__mux4_1 c391 (.A0(net307),
    .A1(net66),
    .A2(net888),
    .A3(net990),
    .S0(net897),
    .S1(net766),
    .X(net308));
 sky130_fd_sc_hd__mux4_2 c392 (.A0(net58),
    .A1(net52),
    .A2(net825),
    .A3(net954),
    .S0(net271),
    .S1(net766),
    .X(net309));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net308),
    .A1(net306),
    .A2(net66),
    .A3(net975),
    .S0(net953),
    .S1(net1022),
    .X(net310));
 sky130_fd_sc_hd__mux4_1 c394 (.A0(net293),
    .A1(net1020),
    .A2(net856),
    .A3(net919),
    .S0(net975),
    .S1(clknet_1_1__leaf_net744),
    .X(net311));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net292),
    .A1(net310),
    .A2(net37),
    .A3(net975),
    .S0(net748),
    .S1(net765),
    .X(net312));
 sky130_fd_sc_hd__and2_2 c396 (.A(net1011),
    .B(net204),
    .X(net313));
 sky130_fd_sc_hd__and3_4 c397 (.A(net81),
    .B(net205),
    .C(net963),
    .X(net314));
 sky130_fd_sc_hd__a2111o_2 c398 (.A1(net984),
    .A2(net85),
    .B1(net314),
    .C1(net191),
    .D1(net963),
    .X(net315));
 sky130_fd_sc_hd__and2_1 c399 (.A(net313),
    .B(net1004),
    .X(net316));
 sky130_fd_sc_hd__and3_2 c400 (.A(net996),
    .B(net75),
    .C(net192),
    .X(net317));
 sky130_fd_sc_hd__and3_2 c401 (.A(net703),
    .B(net316),
    .C(net965),
    .X(net318));
 sky130_fd_sc_hd__and3_1 c402 (.A(net318),
    .B(net968),
    .C(net967),
    .X(net319));
 sky130_fd_sc_hd__and3_2 c403 (.A(net1008),
    .B(net1022),
    .C(net313),
    .X(net900));
 sky130_fd_sc_hd__a2111o_2 c404 (.A1(net1020),
    .A2(net996),
    .B1(net74),
    .C1(net968),
    .D1(net945),
    .X(net320));
 sky130_fd_sc_hd__and3_4 c405 (.A(net968),
    .B(net318),
    .C(net945),
    .X(net321));
 sky130_fd_sc_hd__a2111o_2 c406 (.A1(net320),
    .A2(net314),
    .B1(net945),
    .C1(net967),
    .D1(net996),
    .X(net322));
 sky130_fd_sc_hd__a2111o_2 c407 (.A1(net1004),
    .A2(net939),
    .B1(net963),
    .C1(net945),
    .D1(net1021),
    .X(net323));
 sky130_fd_sc_hd__and3_4 c408 (.A(net961),
    .B(net321),
    .C(net945),
    .X(net324));
 sky130_fd_sc_hd__mux4_2 c409 (.A0(net315),
    .A1(net209),
    .A2(net321),
    .A3(net322),
    .S0(net819),
    .S1(net945),
    .X(net325));
 sky130_fd_sc_hd__mux4_2 c410 (.A0(net74),
    .A1(net322),
    .A2(net321),
    .A3(net968),
    .S0(net324),
    .S1(net945),
    .X(net326));
 sky130_fd_sc_hd__mux4_2 c411 (.A0(net939),
    .A1(net326),
    .A2(net318),
    .A3(net324),
    .S0(net321),
    .S1(net1011),
    .X(net327));
 sky130_fd_sc_hd__mux4_2 c412 (.A0(net323),
    .A1(net325),
    .A2(net320),
    .A3(net207),
    .S0(net967),
    .S1(net945),
    .X(net328));
 sky130_fd_sc_hd__and3_4 c413 (.A(net327),
    .B(net1005),
    .C(net946),
    .X(net929));
 sky130_fd_sc_hd__mux4_2 c414 (.A0(net321),
    .A1(net929),
    .A2(net314),
    .A3(net328),
    .S0(net196),
    .S1(net967),
    .X(net329));
 sky130_fd_sc_hd__mux4_2 c415 (.A0(net201),
    .A1(net328),
    .A2(net329),
    .A3(net322),
    .S0(net318),
    .S1(net945),
    .X(net330));
 sky130_fd_sc_hd__a2111o_1 c416 (.A1(net329),
    .A2(net206),
    .B1(net945),
    .C1(net996),
    .D1(net328),
    .X(net331));
 sky130_fd_sc_hd__mux4_1 c417 (.A0(net204),
    .A1(net326),
    .A2(net206),
    .A3(net331),
    .S0(net322),
    .S1(net946),
    .X(net332));
 sky130_fd_sc_hd__a2111o_2 c418 (.A1(net75),
    .A2(net836),
    .B1(net313),
    .C1(net165),
    .D1(net327),
    .X(net333));
 sky130_fd_sc_hd__dlymetal6s2s_1 c419 (.A(net663),
    .X(net334));
 sky130_fd_sc_hd__and3_1 c420 (.A(net949),
    .B(net207),
    .C(net963),
    .X(net335));
 sky130_fd_sc_hd__and3_2 c421 (.A(net91),
    .B(net313),
    .C(net984),
    .X(net926));
 sky130_fd_sc_hd__and3_1 c422 (.A(net320),
    .B(net996),
    .C(net222),
    .X(net336));
 sky130_fd_sc_hd__a2111o_2 c423 (.A1(net334),
    .A2(net1024),
    .B1(net213),
    .C1(net1021),
    .D1(net75),
    .X(net337));
 sky130_fd_sc_hd__or4bb_4 c424 (.A(net836),
    .B(net320),
    .C_N(net926),
    .D_N(net998),
    .X(net338));
 sky130_fd_sc_hd__and3_2 c425 (.A(net200),
    .B(net333),
    .C(net99),
    .X(net339));
 sky130_fd_sc_hd__mux4_2 c426 (.A0(net80),
    .A1(net337),
    .A2(net192),
    .A3(net335),
    .S0(net320),
    .S1(net963),
    .X(net340));
 sky130_fd_sc_hd__buf_1 c427 (.A(net663),
    .X(net341));
 sky130_fd_sc_hd__a2111o_2 c428 (.A1(net216),
    .A2(net93),
    .B1(net313),
    .C1(net962),
    .D1(net964),
    .X(net342));
 sky130_fd_sc_hd__a2111o_2 c429 (.A1(net202),
    .A2(net327),
    .B1(net337),
    .C1(net192),
    .D1(net99),
    .X(net343));
 sky130_fd_sc_hd__or4bb_1 c430 (.A(net103),
    .B(net937),
    .C_N(net224),
    .D_N(net341),
    .X(net344));
 sky130_fd_sc_hd__a2111o_4 c431 (.A1(net1020),
    .A2(net937),
    .B1(net103),
    .C1(net338),
    .D1(net341),
    .X(net345));
 sky130_fd_sc_hd__sdfbbn_2 c432 (.CLK_N(clknet_4_2_0_clk),
    .D(net325),
    .RESET_B(net342),
    .SCD(net948),
    .SCE(net338),
    .SET_B(net321),
    .Q(net347),
    .Q_N(net346));
 sky130_fd_sc_hd__and3_1 c433 (.A(net337),
    .B(net347),
    .C(net846),
    .X(net348));
 sky130_fd_sc_hd__a2111o_1 c434 (.A1(net335),
    .A2(net221),
    .B1(net948),
    .C1(net1052),
    .D1(net937),
    .X(net349));
 sky130_fd_sc_hd__a2111o_4 c435 (.A1(net339),
    .A2(net937),
    .B1(net968),
    .C1(net663),
    .D1(net698),
    .X(net350));
 sky130_fd_sc_hd__a2111o_1 c436 (.A1(net853),
    .A2(net348),
    .B1(net336),
    .C1(net937),
    .D1(net663),
    .X(net351));
 sky130_fd_sc_hd__a2111o_1 c437 (.A1(net341),
    .A2(net980),
    .B1(net937),
    .C1(net939),
    .D1(net663),
    .X(net352));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(net338),
    .A1(net348),
    .A2(net946),
    .A3(net346),
    .S0(net937),
    .S1(net337),
    .X(net353));
 sky130_fd_sc_hd__mux4_2 c439 (.A0(net353),
    .A1(net348),
    .A2(net213),
    .A3(net937),
    .S0(net209),
    .S1(net819),
    .X(net354));
 sky130_fd_sc_hd__mux4_1 c440 (.A0(net231),
    .A1(net127),
    .A2(net993),
    .A3(net900),
    .S0(net942),
    .S1(net988),
    .X(net355));
 sky130_fd_sc_hd__mux4_1 c441 (.A0(net355),
    .A1(net125),
    .A2(net820),
    .A3(net999),
    .S0(net842),
    .S1(net1055),
    .X(net356));
 sky130_fd_sc_hd__mux4_1 c442 (.A0(net197),
    .A1(net126),
    .A2(net247),
    .A3(net354),
    .S0(net74),
    .S1(net937),
    .X(net357));
 sky130_fd_sc_hd__mux4_1 c443 (.A0(net127),
    .A1(net219),
    .A2(net325),
    .A3(net236),
    .S0(net209),
    .S1(net231),
    .X(net358));
 sky130_fd_sc_hd__mux4_2 c444 (.A0(net994),
    .A1(net338),
    .A2(net103),
    .A3(net339),
    .S0(net979),
    .S1(net655),
    .X(net359));
 sky130_fd_sc_hd__mux4_2 c445 (.A0(net938),
    .A1(net982),
    .A2(net950),
    .A3(net961),
    .S0(net699),
    .S1(net727),
    .X(net360));
 sky130_fd_sc_hd__mux4_1 c446 (.A0(net99),
    .A1(net126),
    .A2(net227),
    .A3(net350),
    .S0(net345),
    .S1(net727),
    .X(net361));
 sky130_fd_sc_hd__mux4_2 c447 (.A0(net208),
    .A1(net321),
    .A2(net949),
    .A3(net190),
    .S0(net75),
    .S1(net217),
    .X(net890));
 sky130_fd_sc_hd__mux4_1 c448 (.A0(net950),
    .A1(net355),
    .A2(net350),
    .A3(net236),
    .S0(net983),
    .S1(net218),
    .X(net362));
 sky130_fd_sc_hd__mux4_1 c449 (.A0(net358),
    .A1(net343),
    .A2(net926),
    .A3(net350),
    .S0(net890),
    .S1(net222),
    .X(net363));
 sky130_fd_sc_hd__mux4_2 c450 (.A0(net75),
    .A1(net994),
    .A2(net91),
    .A3(net993),
    .S0(net346),
    .S1(net948),
    .X(net364));
 sky130_fd_sc_hd__mux4_1 c451 (.A0(net242),
    .A1(net338),
    .A2(net247),
    .A3(net354),
    .S0(net964),
    .S1(net937),
    .X(net365));
 sky130_fd_sc_hd__mux4_1 c452 (.A0(net939),
    .A1(net889),
    .A2(net365),
    .A3(net988),
    .S0(net730),
    .S1(net770),
    .X(net366));
 sky130_fd_sc_hd__sdfbbp_1 c453 (.CLK(clknet_4_3_0_clk),
    .D(net354),
    .RESET_B(net91),
    .SCD(net342),
    .SCE(net358),
    .SET_B(net730),
    .Q(net368),
    .Q_N(net367));
 sky130_fd_sc_hd__mux4_1 c454 (.A0(net365),
    .A1(net359),
    .A2(net1015),
    .A3(net1002),
    .S0(net730),
    .S1(net987),
    .X(net369));
 sky130_fd_sc_hd__mux4_1 c455 (.A0(net336),
    .A1(net325),
    .A2(net365),
    .A3(net1069),
    .S0(net1072),
    .S1(net1058),
    .X(net370));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(net364),
    .A1(net890),
    .A2(net1006),
    .A3(net222),
    .S0(net994),
    .S1(net1068),
    .X(net371));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(net873),
    .A1(net336),
    .A2(net1021),
    .A3(net371),
    .S0(net1055),
    .S1(net1050),
    .X(net372));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(net246),
    .A1(net0),
    .A2(net371),
    .A3(net994),
    .S0(net654),
    .S1(net1062),
    .X(net373));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net206),
    .A1(net350),
    .A2(net365),
    .A3(net359),
    .S0(net771),
    .S1(net773),
    .X(net374));
 sky130_fd_sc_hd__mux4_2 c460 (.A0(net197),
    .A1(net238),
    .A2(net933),
    .A3(net654),
    .S0(net699),
    .S1(net773),
    .X(net375));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net371),
    .A1(net222),
    .A2(net375),
    .A3(net242),
    .S0(net772),
    .S1(net773),
    .X(net376));
 sky130_fd_sc_hd__mux4_1 c462 (.A0(net822),
    .A1(net190),
    .A2(net1000),
    .A3(net926),
    .S0(net1034),
    .S1(net655),
    .X(net377));
 sky130_fd_sc_hd__mux4_1 c463 (.A0(net377),
    .A1(net938),
    .A2(net268),
    .A3(net891),
    .S0(net247),
    .S1(net774),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 c464 (.A0(net948),
    .A1(net984),
    .A2(net367),
    .A3(net735),
    .S0(net745),
    .S1(net771),
    .X(net379));
 sky130_fd_sc_hd__mux4_1 c465 (.A0(net368),
    .A1(net1034),
    .A2(net239),
    .A3(net940),
    .S0(net359),
    .S1(net966),
    .X(net380));
 sky130_fd_sc_hd__mux4_1 c466 (.A0(net227),
    .A1(net324),
    .A2(net125),
    .A3(net938),
    .S0(net1016),
    .S1(net774),
    .X(net381));
 sky130_fd_sc_hd__mux4_1 c467 (.A0(net131),
    .A1(net938),
    .A2(net979),
    .A3(net824),
    .S0(net989),
    .S1(net767),
    .X(net382));
 sky130_fd_sc_hd__mux4_1 c468 (.A0(net359),
    .A1(net350),
    .A2(net227),
    .A3(net952),
    .S0(net958),
    .S1(net988),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 c469 (.A0(net81),
    .A1(net872),
    .A2(net997),
    .A3(net821),
    .S0(net824),
    .S1(net772),
    .X(net384));
 sky130_fd_sc_hd__mux4_1 c470 (.A0(net870),
    .A1(net378),
    .A2(net23),
    .A3(net267),
    .S0(net0),
    .S1(net984),
    .X(net385));
 sky130_fd_sc_hd__mux4_1 c471 (.A0(net129),
    .A1(net239),
    .A2(net81),
    .A3(net323),
    .S0(net270),
    .S1(net217),
    .X(net386));
 sky130_fd_sc_hd__mux4_1 c472 (.A0(net105),
    .A1(net386),
    .A2(net890),
    .A3(net1000),
    .S0(net684),
    .S1(net697),
    .X(net387));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(net261),
    .A1(net387),
    .A2(net263),
    .A3(net948),
    .S0(net676),
    .S1(clknet_1_1__leaf_net775),
    .X(net388));
 sky130_fd_sc_hd__mux4_1 c474 (.A0(net360),
    .A1(net263),
    .A2(net684),
    .A3(net729),
    .S0(net767),
    .S1(clknet_1_1__leaf_net777),
    .X(net389));
 sky130_fd_sc_hd__mux4_1 c475 (.A0(net131),
    .A1(net948),
    .A2(net270),
    .A3(net828),
    .S0(net988),
    .S1(clknet_1_1__leaf_net777),
    .X(net390));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(net190),
    .A1(net1006),
    .A2(net72),
    .A3(net382),
    .S0(net906),
    .S1(clknet_1_0__leaf_net777),
    .X(net391));
 sky130_fd_sc_hd__mux4_2 c477 (.A0(net938),
    .A1(net961),
    .A2(net841),
    .A3(net1006),
    .S0(net824),
    .S1(net940),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(net321),
    .A1(net327),
    .A2(clknet_1_0__leaf_net389),
    .A3(net343),
    .S0(net116),
    .S1(net103),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(net386),
    .A1(net387),
    .A2(net74),
    .A3(net392),
    .S0(net378),
    .S1(net729),
    .X(net394));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net393),
    .A1(net222),
    .A2(clknet_1_0__leaf_net389),
    .A3(net368),
    .S0(net732),
    .S1(net778),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net384),
    .A1(net382),
    .A2(net360),
    .A3(net210),
    .S0(net392),
    .S1(net779),
    .X(net396));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(net387),
    .A1(net938),
    .A2(net900),
    .A3(net396),
    .S0(net979),
    .S1(net779),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net23),
    .A1(net74),
    .A2(net392),
    .A3(clknet_1_1__leaf_net710),
    .S0(clknet_1_1__leaf_net777),
    .S1(net778),
    .X(net398));
 sky130_fd_sc_hd__mux4_1 c484 (.A0(net279),
    .A1(net837),
    .A2(net849),
    .A3(net884),
    .S0(net1051),
    .S1(net1056),
    .X(net399));
 sky130_fd_sc_hd__mux4_1 c485 (.A0(net382),
    .A1(net360),
    .A2(net116),
    .A3(clknet_1_1__leaf_net398),
    .S0(net270),
    .S1(net767),
    .X(net400));
 sky130_fd_sc_hd__mux4_1 c486 (.A0(net343),
    .A1(net866),
    .A2(net269),
    .A3(net30),
    .S0(net246),
    .S1(net779),
    .X(net401));
 sky130_fd_sc_hd__mux4_1 c487 (.A0(net266),
    .A1(net919),
    .A2(clknet_1_0__leaf_net911),
    .A3(net956),
    .S0(net912),
    .S1(net246),
    .X(net402));
 sky130_fd_sc_hd__mux4_1 c488 (.A0(net333),
    .A1(net116),
    .A2(net343),
    .A3(net1018),
    .S0(net236),
    .S1(net729),
    .X(net403));
 sky130_fd_sc_hd__mux4_1 c489 (.A0(clknet_1_0__leaf_net276),
    .A1(clknet_1_1__leaf_net389),
    .A2(net863),
    .A3(net30),
    .S0(net691),
    .S1(net921),
    .X(net404));
 sky130_fd_sc_hd__mux4_1 c490 (.A0(net218),
    .A1(net10),
    .A2(net345),
    .A3(net266),
    .S0(net343),
    .S1(net987),
    .X(net405));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(net403),
    .A1(net926),
    .A2(net248),
    .A3(net247),
    .S0(net691),
    .S1(net757),
    .X(net406));
 sky130_fd_sc_hd__mux4_1 c492 (.A0(net390),
    .A1(net849),
    .A2(net1006),
    .A3(net923),
    .S0(net997),
    .S1(net782),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(net837),
    .A1(net919),
    .A2(net30),
    .A3(net1022),
    .S0(net861),
    .S1(net675),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(net891),
    .A1(net909),
    .A2(clknet_1_0__leaf_net758),
    .A3(net771),
    .S0(net783),
    .S1(net784),
    .X(net409));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(clknet_1_0__leaf_net281),
    .A1(clknet_1_0__leaf_net276),
    .A2(net125),
    .A3(net73),
    .S0(net1041),
    .S1(net784),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(net284),
    .A1(net266),
    .A2(net942),
    .A3(net116),
    .S0(net724),
    .S1(net767),
    .X(net411));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net116),
    .A1(net1018),
    .A2(net248),
    .A3(net908),
    .S0(net695),
    .S1(net784),
    .X(net412));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(net890),
    .A1(net267),
    .A2(net139),
    .A3(net725),
    .S0(net783),
    .S1(net784),
    .X(net413));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(net30),
    .A1(net955),
    .A2(clknet_1_1__leaf_net398),
    .A3(net723),
    .S0(net757),
    .S1(net784),
    .X(net414));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(net360),
    .A1(net1005),
    .A2(net1028),
    .A3(net725),
    .S0(net780),
    .S1(net784),
    .X(net415));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(net395),
    .A1(net923),
    .A2(net415),
    .A3(net982),
    .S0(net30),
    .S1(net782),
    .X(net416));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(net953),
    .A1(net990),
    .A2(net16),
    .A3(net724),
    .S0(net780),
    .S1(net784),
    .X(net417));
 sky130_fd_sc_hd__mux4_2 c503 (.A0(net125),
    .A1(net417),
    .A2(net918),
    .A3(net15),
    .S0(net36),
    .S1(net782),
    .X(net418));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net414),
    .A1(net904),
    .A2(net942),
    .A3(net1018),
    .S0(net761),
    .S1(net767),
    .X(net419));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(net419),
    .A1(net982),
    .A2(net324),
    .A3(net129),
    .S0(net30),
    .S1(net757),
    .X(net420));
 sky130_fd_sc_hd__mux4_1 c526 (.A0(net350),
    .A1(net992),
    .A2(net894),
    .A3(net908),
    .S0(net920),
    .S1(net784),
    .X(net421));
 sky130_fd_sc_hd__mux4_1 c527 (.A0(net834),
    .A1(net284),
    .A2(net312),
    .A3(net304),
    .S0(net894),
    .S1(clknet_1_1__leaf_net901),
    .X(net422));
 sky130_fd_sc_hd__buf_1 c528 (.A(net690),
    .X(net423));
 sky130_fd_sc_hd__or4bb_1 c529 (.A(net87),
    .B(net331),
    .C_N(net1018),
    .D_N(net999),
    .X(net424));
 sky130_fd_sc_hd__and3_1 c530 (.A(net318),
    .B(net197),
    .C(net929),
    .X(net425));
 sky130_fd_sc_hd__a2111o_4 c531 (.A1(net197),
    .A2(net324),
    .B1(net963),
    .C1(net999),
    .D1(net1021),
    .X(net426));
 sky130_fd_sc_hd__a2111o_4 c532 (.A1(net328),
    .A2(net314),
    .B1(net969),
    .C1(net426),
    .D1(net980),
    .X(net427));
 sky130_fd_sc_hd__or4bb_1 c533 (.A(net323),
    .B(net939),
    .C_N(net68),
    .D_N(net672),
    .X(net428));
 sky130_fd_sc_hd__and3_4 c534 (.A(net427),
    .B(net948),
    .C(net980),
    .X(net429));
 sky130_fd_sc_hd__and3_1 c535 (.A(net85),
    .B(net209),
    .C(net1013),
    .X(net430));
 sky130_fd_sc_hd__or4bb_1 c536 (.A(net425),
    .B(net318),
    .C_N(net939),
    .D_N(net965),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_1 c537 (.A(net690),
    .X(net432));
 sky130_fd_sc_hd__and3_1 c538 (.A(net1015),
    .B(net318),
    .C(net994),
    .X(net433));
 sky130_fd_sc_hd__mux4_2 c539 (.A0(net948),
    .A1(net200),
    .A2(net1008),
    .A3(net425),
    .S0(net192),
    .S1(net426),
    .X(net434));
 sky130_fd_sc_hd__sdfrbp_1 c540 (.CLK(clknet_4_0_0_clk),
    .D(net434),
    .RESET_B(net87),
    .SCD(net433),
    .SCE(net947),
    .Q(net436),
    .Q_N(net435));
 sky130_fd_sc_hd__a2111o_4 c541 (.A1(net430),
    .A2(net1024),
    .B1(net426),
    .C1(net969),
    .D1(net429),
    .X(net437));
 sky130_fd_sc_hd__sdfbbn_2 c542 (.CLK_N(clknet_4_2_0_clk),
    .D(net433),
    .RESET_B(net969),
    .SCD(net423),
    .SCE(net85),
    .SET_B(net434),
    .Q(net915),
    .Q_N(net438));
 sky130_fd_sc_hd__sdfbbn_2 c543 (.CLK_N(clknet_4_0_0_clk),
    .D(net1061),
    .RESET_B(net314),
    .SCD(net435),
    .SCE(net87),
    .SET_B(net434),
    .Q(net907),
    .Q_N(net439));
 sky130_fd_sc_hd__a2111o_1 c544 (.A1(net431),
    .A2(net437),
    .B1(net969),
    .C1(net1059),
    .D1(net439),
    .X(net440));
 sky130_fd_sc_hd__a2111o_1 c545 (.A1(net430),
    .A2(net428),
    .B1(net439),
    .C1(net672),
    .D1(net690),
    .X(net441));
 sky130_fd_sc_hd__mux4_2 c546 (.A0(net436),
    .A1(net432),
    .A2(net907),
    .A3(net192),
    .S0(net437),
    .S1(net689),
    .X(net442));
 sky130_fd_sc_hd__a2111o_1 c547 (.A1(net428),
    .A2(net442),
    .B1(net439),
    .C1(net934),
    .D1(net689),
    .X(net443));
 sky130_fd_sc_hd__mux4_1 c548 (.A0(net322),
    .A1(net427),
    .A2(net907),
    .A3(net438),
    .S0(net442),
    .S1(net672),
    .X(net444));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(net968),
    .A1(net326),
    .A2(net434),
    .A3(net442),
    .S0(net672),
    .S1(net785),
    .X(net445));
 sky130_fd_sc_hd__a2111o_2 c550 (.A1(net89),
    .A2(net352),
    .B1(net76),
    .C1(net429),
    .D1(net988),
    .X(net446));
 sky130_fd_sc_hd__a2111o_1 c551 (.A1(net100),
    .A2(net205),
    .B1(net446),
    .C1(net843),
    .D1(net200),
    .X(net447));
 sky130_fd_sc_hd__a2111o_1 c552 (.A1(net192),
    .A2(net929),
    .B1(net334),
    .C1(net980),
    .D1(net196),
    .X(net448));
 sky130_fd_sc_hd__mux4_1 c553 (.A0(net980),
    .A1(net934),
    .A2(net220),
    .A3(net447),
    .S0(net213),
    .S1(net1013),
    .X(net449));
 sky130_fd_sc_hd__a2111o_2 c554 (.A1(net427),
    .A2(net1001),
    .B1(net988),
    .C1(net698),
    .D1(net986),
    .X(net450));
 sky130_fd_sc_hd__mux4_1 c555 (.A0(net96),
    .A1(net342),
    .A2(net1002),
    .A3(net429),
    .S0(net438),
    .S1(net439),
    .X(net451));
 sky130_fd_sc_hd__sdfbbp_1 c556 (.CLK(clknet_4_2_0_clk),
    .D(net846),
    .RESET_B(net342),
    .SCD(net1008),
    .SCE(net934),
    .SET_B(net929),
    .Q(net453),
    .Q_N(net452));
 sky130_fd_sc_hd__a2111o_2 c557 (.A1(net1024),
    .A2(net423),
    .B1(net209),
    .C1(net190),
    .D1(net986),
    .X(net454));
 sky130_fd_sc_hd__mux4_1 c558 (.A0(net453),
    .A1(net334),
    .A2(net703),
    .A3(net442),
    .S0(net965),
    .S1(net986),
    .X(net455));
 sky130_fd_sc_hd__mux4_2 c559 (.A0(net1021),
    .A1(net429),
    .A2(net932),
    .A3(net452),
    .S0(net441),
    .S1(net986),
    .X(net456));
 sky130_fd_sc_hd__mux4_1 c560 (.A0(net703),
    .A1(net842),
    .A2(net1054),
    .A3(net330),
    .S0(net932),
    .S1(net1067),
    .X(net457));
 sky130_fd_sc_hd__a2111o_4 c561 (.A1(net95),
    .A2(net1015),
    .B1(net1014),
    .C1(net698),
    .D1(net986),
    .X(net458));
 sky130_fd_sc_hd__a2111o_2 c562 (.A1(net423),
    .A2(net209),
    .B1(net1021),
    .C1(net458),
    .D1(net454),
    .X(net459));
 sky130_fd_sc_hd__a2111o_1 c563 (.A1(net456),
    .A2(net339),
    .B1(net458),
    .C1(net423),
    .D1(net789),
    .X(net460));
 sky130_fd_sc_hd__a2111o_2 c564 (.A1(net947),
    .A2(net944),
    .B1(net314),
    .C1(net652),
    .D1(net788),
    .X(net461));
 sky130_fd_sc_hd__sdfbbn_2 c565 (.CLK_N(clknet_4_2_0_clk),
    .D(net447),
    .RESET_B(net461),
    .SCD(net458),
    .SCE(net446),
    .SET_B(net944),
    .Q(net896),
    .Q_N(net462));
 sky130_fd_sc_hd__mux4_2 c566 (.A0(net999),
    .A1(net461),
    .A2(net213),
    .A3(net1024),
    .S0(net988),
    .S1(net986),
    .X(net463));
 sky130_fd_sc_hd__a2111o_2 c567 (.A1(net314),
    .A2(net462),
    .B1(net932),
    .C1(net96),
    .D1(net205),
    .X(net464));
 sky130_fd_sc_hd__sdfbbn_1 c568 (.CLK_N(clknet_4_3_0_clk),
    .D(net215),
    .RESET_B(net456),
    .SCD(net460),
    .SCE(net939),
    .SET_B(net651),
    .Q(net466),
    .Q_N(net465));
 sky130_fd_sc_hd__a2111o_1 c569 (.A1(net464),
    .A2(net852),
    .B1(net466),
    .C1(net842),
    .D1(net788),
    .X(net467));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net213),
    .A1(net76),
    .A2(net454),
    .A3(net997),
    .S0(net461),
    .S1(net467),
    .X(net468));
 sky130_fd_sc_hd__mux4_1 c571 (.A0(net467),
    .A1(net429),
    .A2(net932),
    .A3(net464),
    .S0(net652),
    .S1(net790),
    .X(net469));
 sky130_fd_sc_hd__mux4_2 c572 (.A0(net375),
    .A1(net872),
    .A2(net427),
    .A3(net843),
    .S0(net684),
    .S1(net774),
    .X(net470));
 sky130_fd_sc_hd__mux4_2 c573 (.A0(net209),
    .A1(net456),
    .A2(net191),
    .A3(net458),
    .S0(net773),
    .S1(net774),
    .X(net471));
 sky130_fd_sc_hd__mux4_1 c574 (.A0(net442),
    .A1(net110),
    .A2(net345),
    .A3(net364),
    .S0(net962),
    .S1(net684),
    .X(net472));
 sky130_fd_sc_hd__mux4_1 c575 (.A0(net467),
    .A1(net873),
    .A2(net110),
    .A3(net950),
    .S0(net442),
    .S1(net773),
    .X(net473));
 sky130_fd_sc_hd__mux4_1 c576 (.A0(net342),
    .A1(net961),
    .A2(net442),
    .A3(net427),
    .S0(net338),
    .S1(net985),
    .X(net474));
 sky130_fd_sc_hd__mux4_1 c577 (.A0(net1008),
    .A1(net330),
    .A2(net460),
    .A3(net438),
    .S0(net793),
    .S1(net985),
    .X(net475));
 sky130_fd_sc_hd__mux4_2 c578 (.A0(net354),
    .A1(net459),
    .A2(net191),
    .A3(net209),
    .S0(net698),
    .S1(net793),
    .X(net476));
 sky130_fd_sc_hd__mux4_2 c579 (.A0(net863),
    .A1(net907),
    .A2(net967),
    .A3(net941),
    .S0(net944),
    .S1(net985),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c580 (.A0(net873),
    .A1(net470),
    .A2(net426),
    .A3(net364),
    .S0(net932),
    .S1(net698),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c581 (.A0(net339),
    .A1(net948),
    .A2(net330),
    .A3(net477),
    .S0(net238),
    .S1(net795),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(net869),
    .A1(net477),
    .A2(net375),
    .A3(net107),
    .S0(net684),
    .S1(net878),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c583 (.A0(net480),
    .A1(net476),
    .A2(net110),
    .A3(net98),
    .S0(net944),
    .S1(net477),
    .X(net481));
 sky130_fd_sc_hd__mux4_2 c584 (.A0(net330),
    .A1(net465),
    .A2(net375),
    .A3(net999),
    .S0(net698),
    .S1(net773),
    .X(net482));
 sky130_fd_sc_hd__mux4_2 c585 (.A0(net873),
    .A1(net364),
    .A2(net315),
    .A3(net196),
    .S0(net932),
    .S1(net793),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c586 (.A0(net454),
    .A1(net241),
    .A2(net476),
    .A3(net375),
    .S0(net1020),
    .S1(clknet_1_0__leaf_net744),
    .X(net484));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(net460),
    .A1(net448),
    .A2(net364),
    .A3(net477),
    .S0(net98),
    .S1(net985),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c588 (.A0(net217),
    .A1(net869),
    .A2(net126),
    .A3(net929),
    .S0(net878),
    .S1(net793),
    .X(net486));
 sky130_fd_sc_hd__mux4_1 c589 (.A0(net983),
    .A1(net442),
    .A2(net476),
    .A3(net338),
    .S0(net895),
    .S1(net786),
    .X(net487));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(net1011),
    .A1(net426),
    .A2(net460),
    .A3(net941),
    .S0(net960),
    .S1(net985),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(net426),
    .A1(net476),
    .A2(net480),
    .A3(net324),
    .S0(net773),
    .S1(net793),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c592 (.A0(net426),
    .A1(net323),
    .A2(net477),
    .A3(net458),
    .S0(net699),
    .S1(net793),
    .X(net490));
 sky130_fd_sc_hd__mux4_2 c593 (.A0(net454),
    .A1(net490),
    .A2(net477),
    .A3(net941),
    .S0(net932),
    .S1(net686),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c594 (.A0(net205),
    .A1(net217),
    .A2(net268),
    .A3(net931),
    .S0(net989),
    .S1(net732),
    .X(net492));
 sky130_fd_sc_hd__mux4_1 c595 (.A0(net217),
    .A1(net961),
    .A2(net994),
    .A3(net891),
    .S0(net346),
    .S1(net985),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c596 (.A0(net931),
    .A1(net935),
    .A2(net427),
    .A3(net907),
    .S0(net738),
    .S1(net790),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c597 (.A0(net313),
    .A1(net959),
    .A2(net217),
    .A3(net1019),
    .S0(net735),
    .S1(clknet_1_1__leaf_net797),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c598 (.A0(net323),
    .A1(net248),
    .A2(net324),
    .A3(net714),
    .S0(net985),
    .S1(clknet_1_1__leaf_net797),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c599 (.A0(net261),
    .A1(net464),
    .A2(net313),
    .A3(net906),
    .S0(net217),
    .S1(clknet_1_1__leaf_net797),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c600 (.A0(net379),
    .A1(net1025),
    .A2(net931),
    .A3(net263),
    .S0(net239),
    .S1(net1022),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c601 (.A0(net470),
    .A1(net984),
    .A2(net315),
    .A3(net907),
    .S0(net739),
    .S1(clknet_1_1__leaf_net797),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(net196),
    .A1(net364),
    .A2(net462),
    .A3(net1015),
    .S0(net1001),
    .S1(net72),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(net268),
    .A1(net1016),
    .A2(net888),
    .A3(clknet_1_1__leaf_net495),
    .S0(net772),
    .S1(clknet_1_1__leaf_net797),
    .X(net928));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(clknet_1_0__leaf_net495),
    .A1(net843),
    .A2(net1019),
    .A3(net993),
    .S0(clknet_1_0__leaf_net710),
    .S1(net793),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net466),
    .A1(net867),
    .A2(net268),
    .A3(clknet_1_1__leaf_net495),
    .S0(net890),
    .S1(net427),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net1016),
    .A1(net458),
    .A2(clknet_1_1__leaf_net391),
    .A3(net852),
    .S0(net1002),
    .S1(net787),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(net477),
    .A1(clknet_1_0__leaf_net502),
    .A2(net915),
    .A3(net1011),
    .S0(net315),
    .S1(net772),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net863),
    .A1(net68),
    .A2(net941),
    .A3(clknet_1_1__leaf_net502),
    .S0(net737),
    .S1(clknet_1_0__leaf_net777),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c609 (.A0(clknet_1_0__leaf_net502),
    .A1(net944),
    .A2(net872),
    .A3(net346),
    .S0(net741),
    .S1(net986),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c610 (.A0(net396),
    .A1(net315),
    .A2(clknet_1_1__leaf_net502),
    .A3(net940),
    .S0(net961),
    .S1(clknet_1_1__leaf_net798),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net503),
    .A1(clknet_1_1__leaf_net502),
    .A2(clknet_1_1__leaf_net710),
    .A3(clknet_1_1__leaf_net776),
    .S0(clknet_1_1__leaf_net797),
    .S1(clknet_1_1__leaf_net798),
    .X(net508));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(net207),
    .A1(clknet_1_0__leaf_net391),
    .A2(clknet_1_1__leaf_net502),
    .A3(net989),
    .S0(net794),
    .S1(clknet_1_1__leaf_net798),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(net427),
    .A1(clknet_1_0__leaf_net502),
    .A2(net1016),
    .A3(clknet_1_0__leaf_net776),
    .S0(net787),
    .S1(clknet_1_0__leaf_net798),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(net852),
    .A1(clknet_1_0__leaf_net495),
    .A2(net347),
    .A3(net743),
    .S0(clknet_1_0__leaf_net797),
    .S1(clknet_1_0__leaf_net798),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net379),
    .A1(clknet_1_1__leaf_net511),
    .A2(net842),
    .A3(net878),
    .S0(net741),
    .S1(clknet_1_0__leaf_net798),
    .X(net512));
 sky130_fd_sc_hd__mux4_1 c616 (.A0(net199),
    .A1(net863),
    .A2(net267),
    .A3(net890),
    .S0(net728),
    .S1(clknet_1_1__leaf_net879),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(net345),
    .A1(net983),
    .A2(net413),
    .A3(net846),
    .S0(net392),
    .S1(net267),
    .X(net514));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(net324),
    .A1(net190),
    .A2(net247),
    .A3(net843),
    .S0(net1043),
    .S1(net1017),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c619 (.A0(net248),
    .A1(clknet_1_0__leaf_net420),
    .A2(net955),
    .A3(net459),
    .S0(net831),
    .S1(net774),
    .X(net516));
 sky130_fd_sc_hd__mux4_2 c62 (.A0(net867),
    .A1(net858),
    .A2(net849),
    .A3(net869),
    .S0(net832),
    .S1(net865),
    .X(net0));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net68),
    .A1(net1042),
    .A2(net26),
    .A3(net101),
    .S0(net723),
    .S1(net774),
    .X(net517));
 sky130_fd_sc_hd__mux4_2 c621 (.A0(net863),
    .A1(net68),
    .A2(net1014),
    .A3(net154),
    .S0(net932),
    .S1(net728),
    .X(net518));
 sky130_fd_sc_hd__mux4_2 c622 (.A0(net944),
    .A1(net16),
    .A2(net236),
    .A3(net1022),
    .S0(net739),
    .S1(net756),
    .X(net519));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(net405),
    .A1(net413),
    .A2(net459),
    .A3(net82),
    .S0(net955),
    .S1(net1064),
    .X(net520));
 sky130_fd_sc_hd__mux4_2 c624 (.A0(net408),
    .A1(net955),
    .A2(net190),
    .A3(net891),
    .S0(net26),
    .S1(net987),
    .X(net521));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net843),
    .A1(net1030),
    .A2(net270),
    .A3(net931),
    .S0(net743),
    .S1(net795),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net415),
    .A1(net26),
    .A2(net518),
    .A3(net327),
    .S0(net781),
    .S1(net800),
    .X(net523));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(clknet_1_1__leaf_net420),
    .A1(net8),
    .A2(net1084),
    .A3(net154),
    .S0(net742),
    .S1(net783),
    .X(net524));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net459),
    .A1(net493),
    .A2(net458),
    .A3(net993),
    .S0(net781),
    .S1(net793),
    .X(net525));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(net26),
    .A1(net518),
    .A2(net1011),
    .A3(net875),
    .S0(net678),
    .S1(net1047),
    .X(net526));
 sky130_fd_sc_hd__mux4_2 c63 (.A0(net869),
    .A1(net867),
    .A2(net859),
    .A3(net864),
    .S0(net862),
    .S1(net868),
    .X(net922));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net500),
    .A1(net846),
    .A2(net983),
    .A3(net345),
    .S0(net1013),
    .S1(net867),
    .X(net527));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net518),
    .A1(net525),
    .A2(net979),
    .A3(net997),
    .S0(net519),
    .S1(net1075),
    .X(net528));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net236),
    .A1(net875),
    .A2(net471),
    .A3(net517),
    .S0(net518),
    .S1(net728),
    .X(net529));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(net471),
    .A1(net392),
    .A2(net525),
    .A3(net982),
    .S0(net740),
    .S1(net780),
    .X(net530));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net1013),
    .A1(net1030),
    .A2(net728),
    .A3(net740),
    .S0(clknet_1_1__leaf_net744),
    .S1(net781),
    .X(net531));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net531),
    .A1(net896),
    .A2(net1000),
    .A3(net68),
    .S0(net889),
    .S1(net783),
    .X(net532));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net327),
    .A1(net1014),
    .A2(clknet_1_0__leaf_net532),
    .A3(net519),
    .S0(net935),
    .S1(net738),
    .X(net533));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net515),
    .A1(net483),
    .A2(clknet_1_1__leaf_net532),
    .A3(net26),
    .S0(net960),
    .S1(net893),
    .X(net534));
 sky130_fd_sc_hd__mux4_2 c64 (.A0(net862),
    .A1(net860),
    .A2(net840),
    .A3(net871),
    .S0(net990),
    .S1(net858),
    .X(net1));
 sky130_fd_sc_hd__mux4_2 c65 (.A0(net832),
    .A1(net824),
    .A2(net852),
    .A3(net833),
    .S0(net995),
    .S1(net830),
    .X(net2));
 sky130_fd_sc_hd__and2_1 c66 (.A(net831),
    .B(net0),
    .X(net3));
 sky130_fd_sc_hd__or4bb_1 c660 (.A(net1004),
    .B(net437),
    .C_N(net965),
    .D_N(net947),
    .X(net535));
 sky130_fd_sc_hd__or4bb_1 c661 (.A(net947),
    .B(net80),
    .C_N(net1018),
    .D_N(net785),
    .X(net536));
 sky130_fd_sc_hd__or4bb_1 c662 (.A(net80),
    .B(net437),
    .C_N(net929),
    .D_N(net965),
    .X(net537));
 sky130_fd_sc_hd__a2111o_4 c663 (.A1(net1020),
    .A2(net934),
    .B1(net929),
    .C1(net978),
    .D1(net965),
    .X(net538));
 sky130_fd_sc_hd__mux4_2 c664 (.A0(net200),
    .A1(net907),
    .A2(net437),
    .A3(net968),
    .S0(net538),
    .S1(net999),
    .X(net539));
 sky130_fd_sc_hd__or4bb_1 c665 (.A(net1003),
    .B(net537),
    .C_N(net538),
    .D_N(net965),
    .X(net540));
 sky130_fd_sc_hd__a2111o_2 c666 (.A1(net939),
    .A2(net978),
    .B1(net538),
    .C1(net785),
    .D1(net786),
    .X(net882));
 sky130_fd_sc_hd__a2111o_1 c667 (.A1(net191),
    .A2(net1002),
    .B1(net80),
    .C1(net538),
    .D1(net1021),
    .X(net541));
 sky130_fd_sc_hd__sdfrbp_1 c668 (.CLK(clknet_4_0_0_clk),
    .D(net965),
    .RESET_B(net535),
    .SCD(net537),
    .SCE(net929),
    .Q(net543),
    .Q_N(net542));
 sky130_fd_sc_hd__or4bb_1 c669 (.A(net329),
    .B(net535),
    .C_N(net439),
    .D_N(net999),
    .X(net544));
 sky130_fd_sc_hd__and3_1 c67 (.A(net825),
    .B(net821),
    .C(net1013),
    .X(net4));
 sky130_fd_sc_hd__sdfbbp_1 c670 (.CLK(clknet_4_0_0_clk),
    .D(net537),
    .RESET_B(net882),
    .SCD(net437),
    .SCE(net538),
    .SET_B(net785),
    .Q(net546),
    .Q_N(net545));
 sky130_fd_sc_hd__or4bb_4 c671 (.A(net436),
    .B(net439),
    .C_N(net978),
    .D_N(net667),
    .X(net547));
 sky130_fd_sc_hd__or4bb_2 c672 (.A(net997),
    .B(net200),
    .C_N(net978),
    .D_N(net667),
    .X(net548));
 sky130_fd_sc_hd__a2111o_2 c673 (.A1(net68),
    .A2(net200),
    .B1(net548),
    .C1(net934),
    .D1(net439),
    .X(net549));
 sky130_fd_sc_hd__sdfbbn_1 c674 (.CLK_N(clknet_4_0_0_clk),
    .D(net535),
    .RESET_B(net548),
    .SCD(net549),
    .SCE(net965),
    .SET_B(net545),
    .Q(net551),
    .Q_N(net550));
 sky130_fd_sc_hd__a2111o_2 c675 (.A1(net1004),
    .A2(net550),
    .B1(net548),
    .C1(net200),
    .D1(net667),
    .X(net552));
 sky130_fd_sc_hd__a2111o_2 c676 (.A1(net552),
    .A2(net545),
    .B1(net550),
    .C1(net968),
    .D1(net547),
    .X(net553));
 sky130_fd_sc_hd__mux4_2 c677 (.A0(net548),
    .A1(net538),
    .A2(net76),
    .A3(net536),
    .S0(net542),
    .S1(net553),
    .X(net554));
 sky130_fd_sc_hd__mux4_1 c678 (.A0(net543),
    .A1(net554),
    .A2(net536),
    .A3(net316),
    .S0(net551),
    .S1(net552),
    .X(net555));
 sky130_fd_sc_hd__mux4_1 c679 (.A0(net316),
    .A1(net539),
    .A2(net552),
    .A3(net934),
    .S0(net554),
    .S1(net802),
    .X(net556));
 sky130_fd_sc_hd__and2_0 c68 (.A(net864),
    .B(net856),
    .X(net5));
 sky130_fd_sc_hd__mux4_2 c680 (.A0(net551),
    .A1(net548),
    .A2(net552),
    .A3(net538),
    .S0(net667),
    .S1(net801),
    .X(net557));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(net554),
    .A1(net316),
    .A2(net557),
    .A3(net553),
    .S0(net802),
    .S1(net803),
    .X(net558));
 sky130_fd_sc_hd__mux4_1 c682 (.A0(net429),
    .A1(net552),
    .A2(net934),
    .A3(net554),
    .S0(net969),
    .S1(net1008),
    .X(net559));
 sky130_fd_sc_hd__mux4_2 c683 (.A0(net76),
    .A1(net464),
    .A2(net352),
    .A3(net831),
    .S0(net1014),
    .S1(net801),
    .X(net560));
 sky130_fd_sc_hd__mux4_1 c684 (.A0(net950),
    .A1(net554),
    .A2(net352),
    .A3(net446),
    .S0(net429),
    .S1(net801),
    .X(net561));
 sky130_fd_sc_hd__mux4_1 c685 (.A0(net560),
    .A1(net538),
    .A2(net438),
    .A3(net549),
    .S0(net785),
    .S1(net1060),
    .X(net562));
 sky130_fd_sc_hd__mux4_1 c686 (.A0(net541),
    .A1(net1002),
    .A2(net554),
    .A3(net786),
    .S0(net807),
    .S1(net808),
    .X(net563));
 sky130_fd_sc_hd__mux4_2 c687 (.A0(net552),
    .A1(net844),
    .A2(net934),
    .A3(net845),
    .S0(net1005),
    .S1(net808),
    .X(net564));
 sky130_fd_sc_hd__mux4_1 c688 (.A0(net1088),
    .A1(net564),
    .A2(net438),
    .A3(net541),
    .S0(net993),
    .S1(net809),
    .X(net565));
 sky130_fd_sc_hd__mux4_1 c689 (.A0(net348),
    .A1(net554),
    .A2(net437),
    .A3(net994),
    .S0(net439),
    .S1(net806),
    .X(net566));
 sky130_fd_sc_hd__and2_2 c69 (.A(net859),
    .B(net854),
    .X(net6));
 sky130_fd_sc_hd__mux4_2 c690 (.A0(net934),
    .A1(net542),
    .A2(net547),
    .A3(net1017),
    .S0(net786),
    .S1(net792),
    .X(net567));
 sky130_fd_sc_hd__mux4_1 c691 (.A0(net216),
    .A1(net1018),
    .A2(net788),
    .A3(net805),
    .S0(net806),
    .S1(net808),
    .X(net568));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(net329),
    .A1(net541),
    .A2(net461),
    .A3(net939),
    .S0(net554),
    .S1(net1053),
    .X(net569));
 sky130_fd_sc_hd__mux4_1 c693 (.A0(net1008),
    .A1(net568),
    .A2(net554),
    .A3(net1017),
    .S0(net80),
    .S1(net681),
    .X(net570));
 sky130_fd_sc_hd__mux4_2 c694 (.A0(net352),
    .A1(net845),
    .A2(net348),
    .A3(net934),
    .S0(net429),
    .S1(net808),
    .X(net571));
 sky130_fd_sc_hd__mux4_2 c695 (.A0(net543),
    .A1(net329),
    .A2(net107),
    .A3(net571),
    .S0(net694),
    .S1(net801),
    .X(net883));
 sky130_fd_sc_hd__mux4_2 c696 (.A0(net334),
    .A1(net947),
    .A2(net1004),
    .A3(net978),
    .S0(net845),
    .S1(net805),
    .X(net572));
 sky130_fd_sc_hd__mux4_1 c697 (.A0(net446),
    .A1(net841),
    .A2(net557),
    .A3(net883),
    .S0(net694),
    .S1(net1063),
    .X(net573));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(net553),
    .A1(net883),
    .A2(net978),
    .A3(net681),
    .S0(net809),
    .S1(net812),
    .X(net574));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(net461),
    .A1(net571),
    .A2(net536),
    .A3(net568),
    .S0(net553),
    .S1(net805),
    .X(net575));
 sky130_fd_sc_hd__and3_1 c70 (.A(net877),
    .B(net4),
    .C(net859),
    .X(net7));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net224),
    .A1(net883),
    .A2(net76),
    .A3(net554),
    .S0(net813),
    .S1(net814),
    .X(net576));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(net536),
    .A1(net571),
    .A2(clknet_1_0__leaf_net711),
    .A3(net791),
    .S0(net806),
    .S1(net814),
    .X(net577));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net572),
    .A1(clknet_1_0__leaf_net577),
    .A2(net553),
    .A3(net883),
    .S0(net698),
    .S1(net814),
    .X(net578));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(clknet_1_0__leaf_net577),
    .A1(net541),
    .A2(net693),
    .A3(net810),
    .S0(net814),
    .S1(net815),
    .X(net579));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net1004),
    .A1(net242),
    .A2(net567),
    .A3(net572),
    .S0(net950),
    .S1(net681),
    .X(net580));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(net867),
    .A1(net939),
    .A2(net693),
    .A3(net986),
    .S0(clknet_1_0__leaf_net796),
    .S1(net801),
    .X(net581));
 sky130_fd_sc_hd__mux4_1 c706 (.A0(net538),
    .A1(net1003),
    .A2(net936),
    .A3(net947),
    .S0(net883),
    .S1(net458),
    .X(net582));
 sky130_fd_sc_hd__mux4_2 c707 (.A0(net1088),
    .A1(net107),
    .A2(net247),
    .A3(net786),
    .S0(net985),
    .S1(net807),
    .X(net583));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(net996),
    .A1(net965),
    .A2(net107),
    .A3(net547),
    .S0(net768),
    .S1(net804),
    .X(net584));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(net1089),
    .A1(net437),
    .A2(net463),
    .A3(net1005),
    .S0(clknet_1_0__leaf_net711),
    .S1(net986),
    .X(net585));
 sky130_fd_sc_hd__and2_2 c71 (.A(net821),
    .B(net1016),
    .X(net8));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net0),
    .A1(net1012),
    .A2(net547),
    .A3(net583),
    .S0(net126),
    .S1(clknet_1_0__leaf_net744),
    .X(net586));
 sky130_fd_sc_hd__mux4_2 c711 (.A0(net110),
    .A1(net491),
    .A2(net584),
    .A3(net242),
    .S0(net962),
    .S1(net437),
    .X(net587));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net557),
    .A1(net110),
    .A2(net448),
    .A3(net126),
    .S0(net191),
    .S1(net807),
    .X(net588));
 sky130_fd_sc_hd__mux4_1 c713 (.A0(net572),
    .A1(net491),
    .A2(net587),
    .A3(net895),
    .S0(net750),
    .S1(net768),
    .X(net589));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(net338),
    .A1(net241),
    .A2(net882),
    .A3(net978),
    .S0(clknet_1_1__leaf_net577),
    .S1(net804),
    .X(net590));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net437),
    .A1(net1012),
    .A2(net1088),
    .A3(net996),
    .S0(net567),
    .S1(net816),
    .X(net591));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net587),
    .A1(net994),
    .A2(net463),
    .A3(net583),
    .S0(net564),
    .S1(net772),
    .X(net592));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net571),
    .A1(net567),
    .A2(net587),
    .A3(net1008),
    .S0(net786),
    .S1(net788),
    .X(net593));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(net126),
    .A1(net587),
    .A2(net968),
    .A3(net786),
    .S0(clknet_1_1__leaf_net796),
    .S1(net816),
    .X(net594));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net1005),
    .A1(net845),
    .A2(net239),
    .A3(net572),
    .S0(net107),
    .S1(clknet_1_1__leaf_net775),
    .X(net595));
 sky130_fd_sc_hd__and3_4 c72 (.A(net1),
    .B(net860),
    .C(net0),
    .X(net9));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net585),
    .A1(net347),
    .A2(net0),
    .A3(net491),
    .S0(net786),
    .S1(clknet_1_0__leaf_net817),
    .X(net596));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net448),
    .A1(net580),
    .A2(net347),
    .A3(net583),
    .S0(net587),
    .S1(net806),
    .X(net597));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net567),
    .A1(net338),
    .A2(net557),
    .A3(net979),
    .S1(net746),
    .X(net598));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net984),
    .A1(net587),
    .A2(net1071),
    .A3(net1066),
    .S0(net807),
    .S1(net1048),
    .X(net599));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net491),
    .A1(net895),
    .A2(net747),
    .A3(net750),
    .S0(net815),
    .S1(clknet_1_0__leaf_net817),
    .X(net600));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net241),
    .A1(net546),
    .A2(net950),
    .A3(clknet_1_0__leaf_net600),
    .S0(net715),
    .S1(net813),
    .X(net601));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net15),
    .A1(net966),
    .A2(net0),
    .A3(net750),
    .S0(clknet_1_0__leaf_net797),
    .S1(net802),
    .X(net602));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(clknet_1_1__leaf_net577),
    .A1(net931),
    .A2(net219),
    .A3(net560),
    .S0(net882),
    .S1(net686),
    .X(net603));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net591),
    .A1(net581),
    .A2(net549),
    .A3(net845),
    .S0(net720),
    .S1(net806),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(net490),
    .A1(net960),
    .A2(net584),
    .A3(net935),
    .S0(clknet_1_1__leaf_net775),
    .S1(clknet_1_0__leaf_net818),
    .X(net605));
 sky130_fd_sc_hd__and2_2 c73 (.A(net834),
    .B(net864),
    .X(net10));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net841),
    .A1(net501),
    .A2(net211),
    .A3(net933),
    .S0(net900),
    .S1(net739),
    .X(net606));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net497),
    .A1(net984),
    .A2(net857),
    .A3(net458),
    .S0(clknet_1_0__leaf_net602),
    .S1(net539),
    .X(net607));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(net549),
    .A1(net547),
    .A2(net736),
    .A3(net746),
    .S0(net985),
    .S1(clknet_1_1__leaf_net817),
    .X(net608));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net994),
    .A1(net1012),
    .A2(net512),
    .A3(net883),
    .S0(net1002),
    .S1(net463),
    .X(net609));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(clknet_1_0__leaf_net398),
    .A1(net989),
    .A2(clknet_1_0__leaf_net710),
    .A3(net716),
    .S0(net736),
    .S1(net802),
    .X(net610));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net936),
    .A1(net933),
    .A2(net326),
    .A3(net961),
    .S0(clknet_1_1__leaf_net711),
    .S1(net985),
    .X(net611));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(net347),
    .A1(net219),
    .A2(net564),
    .A3(net936),
    .S0(clknet_1_0__leaf_net600),
    .S1(net743),
    .X(net612));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net463),
    .A1(clknet_1_0__leaf_net511),
    .A2(net539),
    .A3(net828),
    .S0(net989),
    .S1(clknet_1_0__leaf_net797),
    .X(net613));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net239),
    .A1(net959),
    .A2(net915),
    .A3(net591),
    .S0(net269),
    .S1(net772),
    .X(net614));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(net326),
    .A1(net936),
    .A2(clknet_1_0__leaf_net879),
    .A3(clknet_1_0__leaf_net776),
    .S0(net810),
    .S1(clknet_1_0__leaf_net818),
    .X(net615));
 sky130_fd_sc_hd__and2_1 c74 (.A(net7),
    .B(net858),
    .X(net11));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(net583),
    .A1(net831),
    .A2(net857),
    .A3(net959),
    .S0(net720),
    .S1(net802),
    .X(net616));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(net606),
    .A1(net560),
    .A2(net933),
    .A3(net966),
    .S0(net929),
    .S1(clknet_1_0__leaf_net797),
    .X(net617));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(net546),
    .A1(net857),
    .A2(net931),
    .A3(net583),
    .S0(net886),
    .S1(net806),
    .X(net618));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(clknet_1_1__leaf_net611),
    .A1(clknet_1_1__leaf_net600),
    .A2(clknet_1_0__leaf_net610),
    .A3(net915),
    .S0(clknet_1_0__leaf_net775),
    .S1(clknet_1_1__leaf_net818),
    .X(net619));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(clknet_1_0__leaf_net611),
    .A1(net979),
    .A2(clknet_1_0__leaf_net595),
    .A3(net720),
    .S0(net886),
    .S1(net739),
    .X(net887));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(clknet_1_0__leaf_net615),
    .A1(net0),
    .A2(net583),
    .A3(net845),
    .S0(clknet_1_1__leaf_net879),
    .S1(net806),
    .X(net620));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net549),
    .A1(clknet_1_1__leaf_net615),
    .A2(clknet_1_0__leaf_net511),
    .A3(net716),
    .S0(net720),
    .S1(net738),
    .X(net621));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(net564),
    .A1(net621),
    .A2(net219),
    .A3(net936),
    .S0(net685),
    .S1(net806),
    .X(net622));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net959),
    .A1(net1005),
    .A2(net392),
    .A3(net997),
    .S0(net1000),
    .S1(net844),
    .X(net623));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net458),
    .A1(net623),
    .A2(net826),
    .A3(net935),
    .S0(clknet_1_1__leaf_net711),
    .S1(net715),
    .X(net624));
 sky130_fd_sc_hd__and3_2 c75 (.A(net823),
    .B(net870),
    .C(net852),
    .X(net12));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(net539),
    .A1(net267),
    .A2(net1013),
    .A3(net624),
    .S0(net154),
    .S1(clknet_1_1__leaf_net818),
    .X(net625));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(clknet_1_0__leaf_net595),
    .A1(net831),
    .A2(net513),
    .A3(clknet_1_1__leaf_net608),
    .S0(net521),
    .S1(clknet_1_0__leaf_net775),
    .X(net626));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net263),
    .A1(net211),
    .A2(net1076),
    .A3(net69),
    .S0(net935),
    .S1(net737),
    .X(net627));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(clknet_1_1__leaf_net602),
    .A1(net1026),
    .A2(net1019),
    .A3(clknet_1_0__leaf_net608),
    .S0(net893),
    .S1(net811),
    .X(net628));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net269),
    .A1(net69),
    .A2(net1005),
    .A3(net932),
    .S0(net962),
    .S1(net736),
    .X(net629));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net876),
    .A1(net628),
    .A2(net960),
    .A3(net1030),
    .S0(net737),
    .S1(net756),
    .X(net630));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net932),
    .A1(net940),
    .A2(net931),
    .A3(net979),
    .S0(net722),
    .S1(net743),
    .X(net631));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(clknet_1_1__leaf_net610),
    .A1(net627),
    .A2(net418),
    .A3(net883),
    .S0(clknet_1_0__leaf_net775),
    .S1(net811),
    .X(net632));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net1013),
    .A1(net933),
    .A2(net886),
    .A3(net893),
    .S0(net793),
    .S1(net815),
    .X(net633));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net969),
    .A1(net633),
    .A2(net8),
    .A3(net828),
    .S0(net761),
    .S1(clknet_1_1__leaf_net818),
    .X(net634));
 sky130_fd_sc_hd__and3_4 c76 (.A(net9),
    .B(net1010),
    .C(net6),
    .X(net13));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net418),
    .A1(net15),
    .A2(net392),
    .A3(net450),
    .S0(net737),
    .S1(net987),
    .X(net635));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net635),
    .A1(net867),
    .A2(net527),
    .A3(net634),
    .S0(net968),
    .S1(net940),
    .X(net636));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net247),
    .A1(net1030),
    .A2(net907),
    .A3(net736),
    .S0(net740),
    .S1(net750),
    .X(net637));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(net317),
    .A1(net935),
    .A2(net16),
    .A3(net521),
    .S0(net247),
    .S1(net915),
    .X(net638));
 sky130_fd_sc_hd__mux4_1 c764 (.A0(net400),
    .A1(net979),
    .A2(net605),
    .A3(net68),
    .S0(net15),
    .S1(net966),
    .X(net639));
 sky130_fd_sc_hd__mux4_1 c765 (.A0(net270),
    .A1(net8),
    .A2(clknet_1_0__leaf_net398),
    .A3(net638),
    .S0(clknet_1_1__leaf_net595),
    .S1(net740),
    .X(net640));
 sky130_fd_sc_hd__mux4_1 c766 (.A0(net88),
    .A1(net154),
    .A2(net622),
    .A3(net637),
    .S0(net959),
    .S1(net1005),
    .X(net641));
 sky130_fd_sc_hd__mux4_1 c767 (.A0(net517),
    .A1(net839),
    .A2(clknet_1_0__leaf_net398),
    .A3(net989),
    .S0(net704),
    .S1(net738),
    .X(net642));
 sky130_fd_sc_hd__mux4_1 c768 (.A0(net547),
    .A1(net1019),
    .A2(net519),
    .A3(net639),
    .S0(net642),
    .S1(net742),
    .X(net643));
 sky130_fd_sc_hd__mux4_1 c769 (.A0(net1019),
    .A1(net638),
    .A2(net678),
    .A3(net722),
    .S0(net781),
    .S1(net793),
    .X(net644));
 sky130_fd_sc_hd__and2_1 c77 (.A(net827),
    .B(net10),
    .X(net14));
 sky130_fd_sc_hd__and3_2 c78 (.A(net10),
    .B(net3),
    .C(net9),
    .X(net15));
 sky130_fd_sc_hd__and3_2 c79 (.A(net15),
    .B(net12),
    .C(net875),
    .X(net16));
 sky130_fd_sc_hd__and3_4 c80 (.A(net13),
    .B(net6),
    .C(net866),
    .X(net17));
 sky130_fd_sc_hd__or4bb_4 c81 (.A(net14),
    .B(net871),
    .C_N(net11),
    .D_N(net970),
    .X(net18));
 sky130_fd_sc_hd__mux4_2 c82 (.A0(net12),
    .A1(net18),
    .A2(net852),
    .A3(net864),
    .S0(net10),
    .S1(net970),
    .X(net19));
 sky130_fd_sc_hd__a2111o_4 c83 (.A1(net16),
    .A2(net18),
    .B1(net970),
    .C1(net13),
    .D1(net19),
    .X(net20));
 sky130_fd_sc_hd__mux4_2 c84 (.A0(net20),
    .A1(net856),
    .A2(net970),
    .A3(net8),
    .S0(net12),
    .S1(net857),
    .X(net21));
 sky130_fd_sc_hd__mux4_2 c85 (.A0(net19),
    .A1(net5),
    .A2(net12),
    .A3(net13),
    .S0(net859),
    .S1(net21),
    .X(net22));
 sky130_fd_sc_hd__or4bb_4 c86 (.A(net8),
    .B(net6),
    .C_N(net970),
    .D_N(net951),
    .X(net23));
 sky130_fd_sc_hd__mux4_2 c87 (.A0(net1044),
    .A1(net3),
    .A2(net23),
    .A3(net951),
    .S0(net4),
    .S1(net21),
    .X(net24));
 sky130_fd_sc_hd__and3_4 c88 (.A(net24),
    .B(net13),
    .C(net850),
    .X(net25));
 sky130_fd_sc_hd__and3_4 c89 (.A(net1010),
    .B(net866),
    .C(net972),
    .X(net26));
 sky130_fd_sc_hd__and3_1 c90 (.A(net874),
    .B(net858),
    .C(net839),
    .X(net27));
 sky130_fd_sc_hd__or4bb_1 c91 (.A(net838),
    .B(net854),
    .C_N(net18),
    .D_N(net1007),
    .X(net28));
 sky130_fd_sc_hd__or4bb_4 c92 (.A(net3),
    .B(net839),
    .C_N(net28),
    .D_N(net837),
    .X(net29));
 sky130_fd_sc_hd__and3_2 c93 (.A(net7),
    .B(net828),
    .C(net972),
    .X(net30));
 sky130_fd_sc_hd__and3_4 c94 (.A(net843),
    .B(net2),
    .C(net862),
    .X(net31));
 sky130_fd_sc_hd__and3_1 c95 (.A(net13),
    .B(net867),
    .C(net24),
    .X(net32));
 sky130_fd_sc_hd__and3_1 c96 (.A(net12),
    .B(net30),
    .C(net867),
    .X(net33));
 sky130_fd_sc_hd__and3_1 c97 (.A(net830),
    .B(net857),
    .C(net26),
    .X(net34));
 sky130_fd_sc_hd__and3_2 c98 (.A(net866),
    .B(net11),
    .C(net12),
    .X(net35));
 sky130_fd_sc_hd__and3_4 c99 (.A(net25),
    .B(net4),
    .C(net856),
    .X(net36));
 sky130_fd_sc_hd__a2111o_1 merge790 (.A1(net333),
    .A2(net221),
    .B1(net206),
    .C1(net336),
    .D1(net337),
    .X(net645));
 sky130_fd_sc_hd__mux4_1 merge791 (.A0(net331),
    .A1(net318),
    .A2(net314),
    .A3(net207),
    .S0(net431),
    .S1(net999),
    .X(net646));
 sky130_fd_sc_hd__and2_0 merge792 (.A(net401),
    .B(net411),
    .X(net647));
 sky130_fd_sc_hd__and2_0 merge793 (.A(net380),
    .B(net381),
    .X(net648));
 sky130_fd_sc_hd__and2_0 merge794 (.A(net230),
    .B(net226),
    .X(net649));
 sky130_fd_sc_hd__and2_0 merge795 (.A(net294),
    .B(net296),
    .X(net650));
 sky130_fd_sc_hd__dfrbp_1 merge796 (.CLK(clknet_4_0_0_clk),
    .D(net468),
    .RESET_B(net457),
    .Q(net652),
    .Q_N(net651));
 sky130_fd_sc_hd__and2_0 merge797 (.A(net604),
    .B(net607),
    .X(net653));
 sky130_fd_sc_hd__dfrbp_1 merge798 (.CLK(clknet_4_3_0_clk),
    .D(net357),
    .RESET_B(net372),
    .Q(net655),
    .Q_N(net654));
 sky130_fd_sc_hd__and2_0 merge799 (.A(net484),
    .B(net485),
    .X(net656));
 sky130_fd_sc_hd__and2_1 merge800 (.A(net272),
    .B(net252),
    .X(net657));
 sky130_fd_sc_hd__and2_0 merge801 (.A(net250),
    .B(net243),
    .X(net658));
 sky130_fd_sc_hd__and2_0 merge802 (.A(net592),
    .B(net593),
    .X(net659));
 sky130_fd_sc_hd__and2_0 merge803 (.A(net644),
    .B(net625),
    .X(net660));
 sky130_fd_sc_hd__and2_0 merge804 (.A(net514),
    .B(net520),
    .X(net661));
 sky130_fd_sc_hd__and2_0 merge805 (.A(net286),
    .B(net283),
    .X(net662));
 sky130_fd_sc_hd__dfrtn_1 merge806 (.CLK_N(clknet_4_2_0_clk),
    .D(net645),
    .RESET_B(net349),
    .Q(net663));
 sky130_fd_sc_hd__dfrtp_4 merge807 (.CLK(clknet_4_11_0_clk),
    .D(net148),
    .RESET_B(net146),
    .Q(net664));
 sky130_fd_sc_hd__and2_0 merge808 (.A(net64),
    .B(net63),
    .X(net665));
 sky130_fd_sc_hd__and2_0 merge809 (.A(net159),
    .B(net163),
    .X(net666));
 sky130_fd_sc_hd__dfrtp_1 merge810 (.CLK(clknet_4_0_0_clk),
    .D(net540),
    .RESET_B(net544),
    .Q(net667));
 sky130_fd_sc_hd__and2_4 merge811 (.A(net188),
    .B(net183),
    .X(net668));
 sky130_fd_sc_hd__and2_0 merge812 (.A(net566),
    .B(net578),
    .X(net669));
 sky130_fd_sc_hd__and2_0 merge813 (.A(net421),
    .B(net422),
    .X(net670));
 sky130_fd_sc_hd__and2_0 merge814 (.A(net492),
    .B(net498),
    .X(net671));
 sky130_fd_sc_hd__dfrtp_1 merge815 (.CLK(clknet_4_2_0_clk),
    .D(net424),
    .RESET_B(net443),
    .Q(net672));
 sky130_fd_sc_hd__and2_0 merge816 (.A(net416),
    .B(net311),
    .X(net673));
 sky130_fd_sc_hd__dfsbp_2 merge817 (.CLK(clknet_4_15_0_clk),
    .SET_B(net666),
    .Q(net675),
    .Q_N(net674));
 sky130_fd_sc_hd__dfsbp_2 merge818 (.CLK(clknet_4_9_0_clk),
    .D(net255),
    .SET_B(net229),
    .Q(net677),
    .Q_N(net676));
 sky130_fd_sc_hd__dfstp_1 merge819 (.CLK(clknet_4_7_0_clk),
    .D(net524),
    .SET_B(net643),
    .Q(net678));
 sky130_fd_sc_hd__and2_0 merge820 (.A(net522),
    .B(net309),
    .X(net679));
 sky130_fd_sc_hd__and2_0 merge821 (.A(net303),
    .B(net298),
    .X(net680));
 sky130_fd_sc_hd__dfstp_1 merge822 (.CLK(clknet_4_1_0_clk),
    .D(net579),
    .SET_B(net569),
    .Q(net681));
 sky130_fd_sc_hd__and2_0 merge823 (.A(net487),
    .B(net620),
    .X(net682));
 sky130_fd_sc_hd__and2_0 merge824 (.A(net488),
    .B(net619),
    .X(net683));
 sky130_fd_sc_hd__dfstp_2 merge825 (.CLK(clknet_4_3_0_clk),
    .D(net244),
    .SET_B(net370),
    .Q(net684));
 sky130_fd_sc_hd__dlrbn_1 merge826 (.D(net489),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net683),
    .Q(net686),
    .Q_N(net685));
 sky130_fd_sc_hd__and2_0 merge827 (.A(net660),
    .B(net507),
    .X(net687));
 sky130_fd_sc_hd__and2_0 merge828 (.A(net523),
    .B(net641),
    .X(net688));
 sky130_fd_sc_hd__dlrbn_1 merge829 (.D(net646),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net440),
    .Q(net690),
    .Q_N(net689));
 sky130_fd_sc_hd__dlrbp_1 merge830 (.D(net662),
    .GATE(clknet_4_12_0_clk),
    .RESET_B(net290),
    .Q(net692),
    .Q_N(net691));
 sky130_fd_sc_hd__dlrbp_1 merge831 (.D(net565),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net669),
    .Q(net694),
    .Q_N(net693));
 sky130_fd_sc_hd__dlrtn_1 merge832 (.D(net673),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net647),
    .Q(net908));
 sky130_fd_sc_hd__dlrtn_1 merge833 (.D(net147),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net143),
    .Q(net695));
 sky130_fd_sc_hd__and2_0 merge834 (.A(net305),
    .B(net680),
    .X(net696));
 sky130_fd_sc_hd__dlrtn_1 merge835 (.D(net649),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net228),
    .Q(net697));
 sky130_fd_sc_hd__dlrtp_4 merge836 (.D(net344),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net351),
    .Q(net698));
 sky130_fd_sc_hd__dlrtp_4 merge837 (.D(net237),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net245),
    .Q(net699));
 sky130_fd_sc_hd__and2_0 merge838 (.A(net504),
    .B(net528),
    .X(net700));
 sky130_fd_sc_hd__and2_0 merge839 (.A(net529),
    .B(net640),
    .X(net701));
 sky130_fd_sc_hd__dlrtp_1 merge840 (.D(net668),
    .GATE(clknet_4_14_0_clk),
    .RESET_B(net182),
    .Q(net702));
 sky130_fd_sc_hd__edfxbp_1 merge841 (.CLK(clknet_4_4_0_clk),
    .DE(net659),
    .Q(net704),
    .Q_N(net598));
 sky130_fd_sc_hd__and2_0 merge842 (.A(net530),
    .B(net636),
    .X(net705));
 sky130_fd_sc_hd__edfxtp_1 merge843 (.CLK(clknet_4_14_0_clk),
    .D(net665),
    .DE(net650),
    .Q(net927));
 sky130_fd_sc_hd__and2_0 merge844 (.A(net533),
    .B(net534),
    .X(net706));
 sky130_fd_sc_hd__and2_0 merge845 (.A(net499),
    .B(net510),
    .X(net707));
 sky130_fd_sc_hd__and2_0 merge846 (.A(net508),
    .B(net505),
    .X(net708));
 sky130_fd_sc_hd__sdlclkp_1 merge847 (.CLK(clknet_4_14_0_clk),
    .GATE(net175),
    .GCLK(net709));
 sky130_fd_sc_hd__sdlclkp_2 merge848 (.CLK(clknet_4_12_0_clk),
    .GATE(net397),
    .SCE(net383),
    .GCLK(net710));
 sky130_fd_sc_hd__sdlclkp_4 merge849 (.CLK(clknet_4_1_0_clk),
    .GATE(net574),
    .SCE(net601),
    .GCLK(net711));
 sky130_fd_sc_hd__and2_0 merge850 (.A(net509),
    .B(net632),
    .X(net712));
 sky130_fd_sc_hd__dfrbp_1 merge851 (.CLK(clknet_4_9_0_clk),
    .D(net256),
    .RESET_B(net282),
    .Q(net714),
    .Q_N(net713));
 sky130_fd_sc_hd__dfrbp_1 merge852 (.CLK(clknet_4_4_0_clk),
    .D(net481),
    .RESET_B(net599),
    .Q(net716),
    .Q_N(net715));
 sky130_fd_sc_hd__and2_0 merge853 (.A(net618),
    .B(net609),
    .X(net717));
 sky130_fd_sc_hd__and2_0 merge854 (.A(net617),
    .B(net612),
    .X(net718));
 sky130_fd_sc_hd__and2_0 merge855 (.A(net613),
    .B(net616),
    .X(net719));
 sky130_fd_sc_hd__dfrtn_1 merge856 (.CLK_N(clknet_4_4_0_clk),
    .D(net582),
    .RESET_B(net718),
    .Q(net720));
 sky130_fd_sc_hd__dfrtp_4 merge857 (.CLK(clknet_4_11_0_clk),
    .D(net260),
    .RESET_B(net181),
    .Q(net899));
 sky130_fd_sc_hd__dfrtp_2 merge858 (.CLK(clknet_4_4_0_clk),
    .D(net474),
    .RESET_B(net712),
    .Q(net878));
 sky130_fd_sc_hd__dfrtp_1 merge859 (.CLK(clknet_4_10_0_clk),
    .D(net249),
    .Q(net251));
 sky130_fd_sc_hd__dfsbp_1 merge860 (.CLK(clknet_4_13_0_clk),
    .D(net409),
    .SET_B(net706),
    .Q(net723),
    .Q_N(net722));
 sky130_fd_sc_hd__dfsbp_1 merge861 (.CLK(clknet_4_12_0_clk),
    .D(net412),
    .SET_B(net410),
    .Q(net725),
    .Q_N(net724));
 sky130_fd_sc_hd__dfstp_1 merge862 (.CLK(clknet_4_5_0_clk),
    .D(net719),
    .SET_B(net717),
    .Q(net886));
 sky130_fd_sc_hd__and2_0 merge863 (.A(net631),
    .B(net626),
    .X(net726));
 sky130_fd_sc_hd__dfstp_2 merge864 (.CLK(clknet_4_8_0_clk),
    .D(net658),
    .SET_B(net356),
    .Q(net727));
 sky130_fd_sc_hd__dfstp_2 merge865 (.CLK(clknet_4_13_0_clk),
    .D(net402),
    .SET_B(net399),
    .Q(net728));
 sky130_fd_sc_hd__dlrbn_1 merge866 (.D(net362),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net648),
    .Q(net730),
    .Q_N(net729));
 sky130_fd_sc_hd__dlrbn_1 merge867 (.D(net265),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net273),
    .Q(net732),
    .Q_N(net731));
 sky130_fd_sc_hd__and2_0 merge868 (.A(net630),
    .B(net629),
    .X(net733));
 sky130_fd_sc_hd__dlrbp_1 merge869 (.D(net670),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net277),
    .Q(net930),
    .Q_N(net734));
 sky130_fd_sc_hd__dlrbp_2 merge870 (.D(net657),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net696),
    .Q(net735),
    .Q_N(net897));
 sky130_fd_sc_hd__dlrtn_1 merge871 (.D(net590),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net726),
    .Q(net736));
 sky130_fd_sc_hd__dlrtn_1 merge872 (.D(net671),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net733),
    .Q(net737));
 sky130_fd_sc_hd__dlrtn_2 merge873 (.D(net682),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net701),
    .Q(net738));
 sky130_fd_sc_hd__dlrtp_2 merge874 (.D(net496),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net653),
    .Q(net739));
 sky130_fd_sc_hd__dlrtp_1 merge875 (.D(net656),
    .GATE(clknet_4_6_0_clk),
    .RESET_B(net486),
    .Q(net895));
 sky130_fd_sc_hd__dlrtp_1 merge876 (.D(net705),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net700),
    .Q(net740));
 sky130_fd_sc_hd__edfxbp_1 merge877 (.CLK(clknet_4_7_0_clk),
    .D(net688),
    .DE(net707),
    .Q(net742),
    .Q_N(net741));
 sky130_fd_sc_hd__edfxtp_1 merge878 (.CLK(clknet_4_7_0_clk),
    .D(net687),
    .DE(net708),
    .Q(net743));
 sky130_fd_sc_hd__sdlclkp_1 merge879 (.CLK(clknet_4_5_0_clk),
    .GATE(net479),
    .SCE(net614),
    .GCLK(net879));
 sky130_fd_sc_hd__sdlclkp_2 merge880 (.CLK(clknet_4_7_0_clk),
    .GATE(net679),
    .SCE(net482),
    .GCLK(net744));
 sky130_fd_sc_hd__sdlclkp_4 merge881 (.CLK(clknet_4_10_0_clk),
    .GATE(net234),
    .GCLK(net235));
 sky130_fd_sc_hd__dfrbp_1 merge882 (.CLK(clknet_4_4_0_clk),
    .D(net597),
    .RESET_B(net596),
    .Q(net747),
    .Q_N(net746));
 sky130_fd_sc_hd__dfrbp_2 merge883 (.CLK(clknet_4_15_0_clk),
    .D(net184),
    .RESET_B(net295),
    .Q(net749),
    .Q_N(net748));
 sky130_fd_sc_hd__dfrtn_1 merge884 (.CLK_N(clknet_4_7_0_clk),
    .D(net661),
    .RESET_B(net526),
    .Q(net893));
 sky130_fd_sc_hd__dfrtp_2 merge885 (.CLK(clknet_4_1_0_clk),
    .D(net588),
    .RESET_B(net586),
    .Q(net750));
 sky130_fd_sc_hd__dfxbp_1 s886 (.CLK(clknet_4_11_0_clk),
    .D(net57),
    .Q(net752),
    .Q_N(net751));
 sky130_fd_sc_hd__dfxbp_1 s887 (.CLK(clknet_4_10_0_clk),
    .D(net144),
    .Q(net754),
    .Q_N(net753));
 sky130_fd_sc_hd__dfxtp_1 s888 (.CLK(clknet_4_14_0_clk),
    .D(net153),
    .Q(net755));
 sky130_fd_sc_hd__dfxtp_2 s889 (.CLK(clknet_4_15_0_clk),
    .D(net167),
    .Q(net756));
 sky130_fd_sc_hd__dfxtp_2 s890 (.CLK(clknet_4_15_0_clk),
    .D(net168),
    .Q(net757));
 sky130_fd_sc_hd__dlclkp_1 s891 (.CLK(clknet_4_15_0_clk),
    .GATE(net169),
    .GCLK(net758));
 sky130_fd_sc_hd__dlclkp_2 s892 (.CLK(clknet_4_11_0_clk),
    .GATE(net172),
    .GCLK(net759));
 sky130_fd_sc_hd__dlclkp_4 s893 (.CLK(clknet_4_11_0_clk),
    .GATE(net178),
    .GCLK(net901));
 sky130_fd_sc_hd__dlxbn_2 s894 (.D(net253),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net761),
    .Q_N(net760));
 sky130_fd_sc_hd__dlxbn_1 s895 (.D(net274),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net920),
    .Q_N(net762));
 sky130_fd_sc_hd__dlxbp_1 s896 (.D(net287),
    .GATE(clknet_4_13_0_clk),
    .Q(net925),
    .Q_N(net763));
 sky130_fd_sc_hd__dlxtn_1 s897 (.D(net288),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net764));
 sky130_fd_sc_hd__dlxtn_1 s898 (.D(net291),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net765));
 sky130_fd_sc_hd__dlxtn_1 s899 (.D(net301),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net766));
 sky130_fd_sc_hd__dlxtp_1 s900 (.D(net332),
    .GATE(clknet_4_2_0_clk),
    .Q(net767));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s901 (.D(net361),
    .SLEEP_B(clknet_4_3_0_clk),
    .Q(net768));
 sky130_fd_sc_hd__dfxbp_1 s902 (.CLK(clknet_4_3_0_clk),
    .D(net363),
    .Q(net770),
    .Q_N(net769));
 sky130_fd_sc_hd__dfxbp_1 s903 (.CLK(clknet_4_13_0_clk),
    .D(net366),
    .Q(net921),
    .Q_N(net771));
 sky130_fd_sc_hd__dfxtp_2 s904 (.CLK(clknet_4_6_0_clk),
    .D(net369),
    .Q(net772));
 sky130_fd_sc_hd__dfxtp_2 s905 (.CLK(clknet_4_3_0_clk),
    .D(net373),
    .Q(net773));
 sky130_fd_sc_hd__dfxtp_2 s906 (.CLK(clknet_4_6_0_clk),
    .D(net374),
    .Q(net774));
 sky130_fd_sc_hd__dlclkp_1 s907 (.CLK(clknet_4_6_0_clk),
    .GATE(net376),
    .GCLK(net775));
 sky130_fd_sc_hd__dlclkp_2 s908 (.CLK(clknet_4_6_0_clk),
    .GATE(net385),
    .GCLK(net776));
 sky130_fd_sc_hd__dlclkp_4 s909 (.CLK(clknet_4_12_0_clk),
    .GATE(net388),
    .GCLK(net777));
 sky130_fd_sc_hd__dlxbn_1 s910 (.D(net394),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net779),
    .Q_N(net778));
 sky130_fd_sc_hd__dlxbn_1 s911 (.D(net404),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net781),
    .Q_N(net780));
 sky130_fd_sc_hd__dlxbp_1 s912 (.D(net406),
    .GATE(clknet_4_12_0_clk),
    .Q(net783),
    .Q_N(net782));
 sky130_fd_sc_hd__dlxtn_2 s913 (.D(net407),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net784));
 sky130_fd_sc_hd__dlxtn_1 s914 (.D(net444),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net785));
 sky130_fd_sc_hd__dlxtn_2 s915 (.D(net445),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net786));
 sky130_fd_sc_hd__dlxtp_1 s916 (.D(net449),
    .GATE(clknet_4_2_0_clk),
    .Q(net787));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s917 (.D(net451),
    .SLEEP_B(clknet_4_0_0_clk),
    .Q(net788));
 sky130_fd_sc_hd__dfxbp_1 s918 (.CLK(clknet_4_2_0_clk),
    .D(net455),
    .Q(net790),
    .Q_N(net789));
 sky130_fd_sc_hd__dfxbp_1 s919 (.CLK(clknet_4_0_0_clk),
    .D(net469),
    .Q(net792),
    .Q_N(net791));
 sky130_fd_sc_hd__dfxtp_4 s920 (.CLK(clknet_4_3_0_clk),
    .D(net472),
    .Q(net793));
 sky130_fd_sc_hd__dfxtp_1 s921 (.CLK(clknet_4_1_0_clk),
    .D(net473),
    .Q(net794));
 sky130_fd_sc_hd__dfxtp_1 s922 (.CLK(clknet_4_3_0_clk),
    .D(net475),
    .Q(net795));
 sky130_fd_sc_hd__dlclkp_1 s923 (.CLK(clknet_4_1_0_clk),
    .GATE(net478),
    .GCLK(net796));
 sky130_fd_sc_hd__dlclkp_2 s924 (.CLK(clknet_4_4_0_clk),
    .GATE(net494),
    .GCLK(net797));
 sky130_fd_sc_hd__dlclkp_4 s925 (.CLK(clknet_4_6_0_clk),
    .GATE(net506),
    .GCLK(net798));
 sky130_fd_sc_hd__dlxbn_1 s926 (.D(net516),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net800),
    .Q_N(net799));
 sky130_fd_sc_hd__dlxbn_2 s927 (.D(net555),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net802),
    .Q_N(net801));
 sky130_fd_sc_hd__dlxbp_1 s928 (.D(net556),
    .GATE(clknet_4_0_0_clk),
    .Q(net804),
    .Q_N(net803));
 sky130_fd_sc_hd__dlxtn_1 s929 (.D(net558),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net805));
 sky130_fd_sc_hd__dlxtn_2 s930 (.D(net559),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net806));
 sky130_fd_sc_hd__dlxtn_1 s931 (.D(net561),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net807));
 sky130_fd_sc_hd__dlxtp_1 s932 (.D(net562),
    .GATE(clknet_4_0_0_clk),
    .Q(net808));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s933 (.D(net563),
    .SLEEP_B(clknet_4_1_0_clk),
    .Q(net809));
 sky130_fd_sc_hd__dfxbp_1 s934 (.CLK(clknet_4_5_0_clk),
    .D(net570),
    .Q(net811),
    .Q_N(net810));
 sky130_fd_sc_hd__dfxbp_1 s935 (.CLK(clknet_4_1_0_clk),
    .D(net573),
    .Q(net813),
    .Q_N(net812));
 sky130_fd_sc_hd__dfxtp_1 s936 (.CLK(clknet_4_0_0_clk),
    .D(net575),
    .Q(net814));
 sky130_fd_sc_hd__dfxtp_1 s937 (.CLK(clknet_4_1_0_clk),
    .D(net576),
    .Q(net815));
 sky130_fd_sc_hd__dfxtp_1 s938 (.CLK(clknet_4_4_0_clk),
    .D(net589),
    .Q(net816));
 sky130_fd_sc_hd__dlclkp_1 s939 (.CLK(clknet_4_4_0_clk),
    .GATE(net594),
    .GCLK(net817));
 sky130_fd_sc_hd__dlclkp_2 s940 (.CLK(clknet_4_4_0_clk),
    .GATE(net603),
    .GCLK(net818));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(in0),
    .X(net165));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(in1),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(in10),
    .X(net703));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(in11),
    .X(net819));
 sky130_fd_sc_hd__buf_1 input5 (.A(in12),
    .X(net820));
 sky130_fd_sc_hd__buf_2 input6 (.A(in13),
    .X(net821));
 sky130_fd_sc_hd__buf_1 input7 (.A(in14),
    .X(net822));
 sky130_fd_sc_hd__buf_2 input8 (.A(in15),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(in16),
    .X(net824));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(in17),
    .X(net825));
 sky130_fd_sc_hd__buf_2 input11 (.A(in18),
    .X(net826));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(in19),
    .X(net827));
 sky130_fd_sc_hd__buf_2 input13 (.A(in2),
    .X(net828));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(in20),
    .X(net829));
 sky130_fd_sc_hd__buf_2 input15 (.A(in21),
    .X(net830));
 sky130_fd_sc_hd__buf_4 input16 (.A(in22),
    .X(net831));
 sky130_fd_sc_hd__buf_2 input17 (.A(in23),
    .X(net832));
 sky130_fd_sc_hd__buf_2 input18 (.A(in24),
    .X(net833));
 sky130_fd_sc_hd__buf_4 input19 (.A(in25),
    .X(net834));
 sky130_fd_sc_hd__buf_2 input20 (.A(in26),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(in27),
    .X(net836));
 sky130_fd_sc_hd__buf_4 input22 (.A(in28),
    .X(net837));
 sky130_fd_sc_hd__buf_2 input23 (.A(in29),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(in3),
    .X(net839));
 sky130_fd_sc_hd__buf_2 input25 (.A(in30),
    .X(net840));
 sky130_fd_sc_hd__clkbuf_4 input26 (.A(in31),
    .X(net841));
 sky130_fd_sc_hd__buf_4 input27 (.A(in32),
    .X(net842));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(in33),
    .X(net843));
 sky130_fd_sc_hd__buf_4 input29 (.A(in34),
    .X(net844));
 sky130_fd_sc_hd__clkbuf_4 input30 (.A(in35),
    .X(net845));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(in36),
    .X(net846));
 sky130_fd_sc_hd__buf_2 input32 (.A(in37),
    .X(net847));
 sky130_fd_sc_hd__buf_2 input33 (.A(in38),
    .X(net848));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(in39),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(in4),
    .X(net850));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(in40),
    .X(net851));
 sky130_fd_sc_hd__clkbuf_4 input37 (.A(in41),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(in42),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(in43),
    .X(net854));
 sky130_fd_sc_hd__buf_1 input40 (.A(in44),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_4 input41 (.A(in45),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(in46),
    .X(net857));
 sky130_fd_sc_hd__buf_2 input43 (.A(in47),
    .X(net858));
 sky130_fd_sc_hd__buf_4 input44 (.A(in48),
    .X(net859));
 sky130_fd_sc_hd__dlymetal6s2s_1 input45 (.A(in49),
    .X(net860));
 sky130_fd_sc_hd__buf_2 input46 (.A(in5),
    .X(net861));
 sky130_fd_sc_hd__buf_8 input47 (.A(in50),
    .X(net862));
 sky130_fd_sc_hd__buf_4 input48 (.A(in51),
    .X(net863));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(in52),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_4 input50 (.A(in53),
    .X(net865));
 sky130_fd_sc_hd__buf_2 input51 (.A(in54),
    .X(net866));
 sky130_fd_sc_hd__buf_6 input52 (.A(in55),
    .X(net867));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(in56),
    .X(net868));
 sky130_fd_sc_hd__buf_6 input54 (.A(in57),
    .X(net869));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(in58),
    .X(net870));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(in59),
    .X(net871));
 sky130_fd_sc_hd__buf_2 input57 (.A(in6),
    .X(net872));
 sky130_fd_sc_hd__buf_2 input58 (.A(in60),
    .X(net873));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(in61),
    .X(net874));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(in7),
    .X(net875));
 sky130_fd_sc_hd__buf_2 input61 (.A(in8),
    .X(net876));
 sky130_fd_sc_hd__dlymetal6s2s_1 input62 (.A(in9),
    .X(net877));
 sky130_fd_sc_hd__buf_2 output63 (.A(net878),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(clknet_1_0__leaf_net879),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output65 (.A(net1083),
    .X(out10));
 sky130_fd_sc_hd__clkbuf_4 output66 (.A(net881),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output67 (.A(net882),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output68 (.A(net883),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output69 (.A(net1030),
    .X(out17));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net885),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output71 (.A(net886),
    .X(out19));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net887),
    .X(out2));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net888),
    .X(out20));
 sky130_fd_sc_hd__clkbuf_4 output74 (.A(net889),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output75 (.A(net890),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output76 (.A(net891),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output77 (.A(net942),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output78 (.A(net893),
    .X(out25));
 sky130_fd_sc_hd__buf_2 output79 (.A(net894),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output80 (.A(net895),
    .X(out27));
 sky130_fd_sc_hd__buf_2 output81 (.A(net896),
    .X(out28));
 sky130_fd_sc_hd__clkbuf_4 output82 (.A(net897),
    .X(out29));
 sky130_fd_sc_hd__clkbuf_4 output83 (.A(net898),
    .X(out3));
 sky130_fd_sc_hd__clkbuf_4 output84 (.A(net899),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output85 (.A(net946),
    .X(out31));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(clknet_1_1__leaf_net901),
    .X(out32));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(clknet_1_1__leaf_net902),
    .X(out34));
 sky130_fd_sc_hd__clkbuf_4 output88 (.A(net981),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output89 (.A(net904),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(clknet_1_1__leaf_net905),
    .X(out37));
 sky130_fd_sc_hd__buf_2 output91 (.A(net933),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output92 (.A(net907),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output93 (.A(net908),
    .X(out41));
 sky130_fd_sc_hd__buf_2 output94 (.A(net931),
    .X(out42));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(clknet_1_1__leaf_net910),
    .X(out43));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(clknet_1_1__leaf_net911),
    .X(out44));
 sky130_fd_sc_hd__buf_2 output97 (.A(net912),
    .X(out45));
 sky130_fd_sc_hd__clkbuf_4 output98 (.A(net913),
    .X(out46));
 sky130_fd_sc_hd__clkbuf_4 output99 (.A(net952),
    .X(out48));
 sky130_fd_sc_hd__buf_2 output100 (.A(net915),
    .X(out5));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(net916),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output102 (.A(net917),
    .X(out51));
 sky130_fd_sc_hd__buf_2 output103 (.A(net918),
    .X(out52));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net943),
    .X(out53));
 sky130_fd_sc_hd__buf_2 output105 (.A(net920),
    .X(out54));
 sky130_fd_sc_hd__buf_2 output106 (.A(net921),
    .X(out55));
 sky130_fd_sc_hd__clkbuf_4 output107 (.A(net922),
    .X(out56));
 sky130_fd_sc_hd__buf_2 output108 (.A(net923),
    .X(out57));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(clknet_1_1__leaf_net924),
    .X(out58));
 sky130_fd_sc_hd__buf_2 output110 (.A(net925),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output111 (.A(net926),
    .X(out60));
 sky130_fd_sc_hd__clkbuf_4 output112 (.A(net927),
    .X(out61));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(net928),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output114 (.A(net929),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output115 (.A(net930),
    .X(out9));
 sky130_fd_sc_hd__buf_4 fanout116 (.A(net909),
    .X(net931));
 sky130_fd_sc_hd__buf_4 fanout117 (.A(net450),
    .X(net932));
 sky130_fd_sc_hd__clkbuf_4 fanout118 (.A(net906),
    .X(net933));
 sky130_fd_sc_hd__clkbuf_4 fanout119 (.A(net441),
    .X(net934));
 sky130_fd_sc_hd__buf_4 fanout120 (.A(net122),
    .X(net935));
 sky130_fd_sc_hd__buf_4 fanout121 (.A(net105),
    .X(net936));
 sky130_fd_sc_hd__clkbuf_4 fanout122 (.A(net340),
    .X(net937));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout123 (.A(net340),
    .X(net938));
 sky130_fd_sc_hd__clkbuf_4 fanout124 (.A(net319),
    .X(net939));
 sky130_fd_sc_hd__clkbuf_2 fanout125 (.A(net319),
    .X(net940));
 sky130_fd_sc_hd__clkbuf_4 fanout126 (.A(net942),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_4 fanout127 (.A(net892),
    .X(net942));
 sky130_fd_sc_hd__clkbuf_4 fanout128 (.A(net919),
    .X(net943));
 sky130_fd_sc_hd__buf_4 fanout129 (.A(net212),
    .X(net944));
 sky130_fd_sc_hd__buf_2 fanout130 (.A(net946),
    .X(net945));
 sky130_fd_sc_hd__clkbuf_2 fanout131 (.A(net947),
    .X(net946));
 sky130_fd_sc_hd__buf_2 fanout132 (.A(net900),
    .X(net947));
 sky130_fd_sc_hd__clkbuf_4 fanout133 (.A(net210),
    .X(net948));
 sky130_fd_sc_hd__clkbuf_4 fanout134 (.A(net101),
    .X(net949));
 sky130_fd_sc_hd__clkbuf_4 fanout135 (.A(net220),
    .X(net950));
 sky130_fd_sc_hd__buf_8 fanout136 (.A(net22),
    .X(net951));
 sky130_fd_sc_hd__buf_4 fanout137 (.A(net914),
    .X(net952));
 sky130_fd_sc_hd__clkbuf_2 fanout138 (.A(net914),
    .X(net953));
 sky130_fd_sc_hd__clkbuf_4 fanout139 (.A(net894),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_4 fanout140 (.A(net278),
    .X(net955));
 sky130_fd_sc_hd__clkbuf_2 fanout141 (.A(net278),
    .X(net956));
 sky130_fd_sc_hd__clkbuf_4 fanout142 (.A(net958),
    .X(net957));
 sky130_fd_sc_hd__clkbuf_4 fanout143 (.A(net959),
    .X(net958));
 sky130_fd_sc_hd__buf_2 fanout144 (.A(net137),
    .X(net959));
 sky130_fd_sc_hd__clkbuf_8 fanout145 (.A(net881),
    .X(net960));
 sky130_fd_sc_hd__buf_4 fanout146 (.A(net88),
    .X(net961));
 sky130_fd_sc_hd__buf_4 fanout147 (.A(net211),
    .X(net962));
 sky130_fd_sc_hd__clkbuf_4 fanout148 (.A(net964),
    .X(net963));
 sky130_fd_sc_hd__buf_2 fanout149 (.A(net966),
    .X(net964));
 sky130_fd_sc_hd__clkbuf_4 fanout150 (.A(net966),
    .X(net965));
 sky130_fd_sc_hd__buf_4 fanout151 (.A(net203),
    .X(net966));
 sky130_fd_sc_hd__buf_4 fanout152 (.A(net199),
    .X(net967));
 sky130_fd_sc_hd__buf_4 fanout153 (.A(net317),
    .X(net968));
 sky130_fd_sc_hd__buf_6 fanout154 (.A(net82),
    .X(net969));
 sky130_fd_sc_hd__buf_8 fanout155 (.A(net971),
    .X(net970));
 sky130_fd_sc_hd__buf_8 fanout156 (.A(net17),
    .X(net971));
 sky130_fd_sc_hd__clkbuf_4 fanout157 (.A(net17),
    .X(net972));
 sky130_fd_sc_hd__buf_1 fanout158 (.A(net17),
    .X(net973));
 sky130_fd_sc_hd__buf_4 fanout159 (.A(net195),
    .X(net974));
 sky130_fd_sc_hd__clkbuf_2 fanout160 (.A(net195),
    .X(net975));
 sky130_fd_sc_hd__buf_2 fanout161 (.A(net978),
    .X(net976));
 sky130_fd_sc_hd__clkbuf_2 fanout162 (.A(net978),
    .X(net977));
 sky130_fd_sc_hd__clkbuf_4 fanout163 (.A(net979),
    .X(net978));
 sky130_fd_sc_hd__buf_4 fanout164 (.A(net189),
    .X(net979));
 sky130_fd_sc_hd__clkbuf_4 fanout165 (.A(net77),
    .X(net980));
 sky130_fd_sc_hd__buf_4 fanout166 (.A(net982),
    .X(net981));
 sky130_fd_sc_hd__clkbuf_4 fanout167 (.A(net903),
    .X(net982));
 sky130_fd_sc_hd__buf_4 fanout168 (.A(net73),
    .X(net983));
 sky130_fd_sc_hd__buf_4 fanout169 (.A(net72),
    .X(net984));
 sky130_fd_sc_hd__buf_4 fanout170 (.A(net794),
    .X(net985));
 sky130_fd_sc_hd__clkbuf_4 fanout171 (.A(net787),
    .X(net986));
 sky130_fd_sc_hd__clkbuf_2 max_cap172 (.A(net768),
    .X(net987));
 sky130_fd_sc_hd__clkbuf_8 fanout173 (.A(net697),
    .X(net988));
 sky130_fd_sc_hd__buf_4 fanout174 (.A(net695),
    .X(net989));
 sky130_fd_sc_hd__buf_8 fanout175 (.A(net922),
    .X(net990));
 sky130_fd_sc_hd__clkbuf_4 fanout176 (.A(net70),
    .X(net991));
 sky130_fd_sc_hd__buf_2 fanout177 (.A(net70),
    .X(net992));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(net69),
    .X(net993));
 sky130_fd_sc_hd__buf_4 fanout179 (.A(net824),
    .X(net994));
 sky130_fd_sc_hd__clkbuf_4 fanout180 (.A(net823),
    .X(net995));
 sky130_fd_sc_hd__clkbuf_4 fanout181 (.A(net822),
    .X(net996));
 sky130_fd_sc_hd__clkbuf_8 fanout182 (.A(net877),
    .X(net997));
 sky130_fd_sc_hd__buf_4 fanout183 (.A(net999),
    .X(net998));
 sky130_fd_sc_hd__buf_4 fanout184 (.A(net1000),
    .X(net999));
 sky130_fd_sc_hd__buf_4 fanout185 (.A(net876),
    .X(net1000));
 sky130_fd_sc_hd__clkbuf_4 fanout186 (.A(net875),
    .X(net1001));
 sky130_fd_sc_hd__buf_4 fanout187 (.A(net821),
    .X(net1002));
 sky130_fd_sc_hd__buf_4 fanout188 (.A(net872),
    .X(net1003));
 sky130_fd_sc_hd__clkbuf_4 fanout189 (.A(net820),
    .X(net1004));
 sky130_fd_sc_hd__buf_4 fanout190 (.A(net861),
    .X(net1005));
 sky130_fd_sc_hd__buf_4 fanout191 (.A(net855),
    .X(net1006));
 sky130_fd_sc_hd__buf_2 fanout192 (.A(net855),
    .X(net1007));
 sky130_fd_sc_hd__clkbuf_4 fanout193 (.A(net819),
    .X(net1008));
 sky130_fd_sc_hd__clkbuf_4 fanout194 (.A(net851),
    .X(net1009));
 sky130_fd_sc_hd__clkbuf_2 fanout195 (.A(net851),
    .X(net1010));
 sky130_fd_sc_hd__buf_4 fanout196 (.A(net850),
    .X(net1011));
 sky130_fd_sc_hd__buf_4 fanout197 (.A(net848),
    .X(net1012));
 sky130_fd_sc_hd__buf_4 fanout198 (.A(net839),
    .X(net1013));
 sky130_fd_sc_hd__clkbuf_8 fanout199 (.A(net835),
    .X(net1014));
 sky130_fd_sc_hd__buf_4 fanout200 (.A(net176),
    .X(net1015));
 sky130_fd_sc_hd__clkbuf_2 fanout201 (.A(net176),
    .X(net1016));
 sky130_fd_sc_hd__buf_4 fanout202 (.A(net830),
    .X(net1017));
 sky130_fd_sc_hd__buf_4 fanout203 (.A(net829),
    .X(net1018));
 sky130_fd_sc_hd__clkbuf_2 fanout204 (.A(net829),
    .X(net1019));
 sky130_fd_sc_hd__clkbuf_8 fanout205 (.A(net828),
    .X(net1020));
 sky130_fd_sc_hd__clkbuf_4 fanout206 (.A(net1022),
    .X(net1021));
 sky130_fd_sc_hd__clkbuf_8 fanout207 (.A(net826),
    .X(net1022));
 sky130_fd_sc_hd__buf_4 fanout208 (.A(net825),
    .X(net1023));
 sky130_fd_sc_hd__clkbuf_4 fanout209 (.A(net165),
    .X(net1024));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net818 (.A(net818),
    .X(clknet_0_net818));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net818 (.A(clknet_0_net818),
    .X(clknet_1_0__leaf_net818));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net818 (.A(clknet_0_net818),
    .X(clknet_1_1__leaf_net818));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net615 (.A(net615),
    .X(clknet_0_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net615 (.A(clknet_0_net615),
    .X(clknet_1_0__leaf_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net615 (.A(clknet_0_net615),
    .X(clknet_1_1__leaf_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net817 (.A(net817),
    .X(clknet_0_net817));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net817 (.A(clknet_0_net817),
    .X(clknet_1_0__leaf_net817));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net817 (.A(clknet_0_net817),
    .X(clknet_1_1__leaf_net817));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net608 (.A(net608),
    .X(clknet_0_net608));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net608 (.A(clknet_0_net608),
    .X(clknet_1_0__leaf_net608));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net608 (.A(clknet_0_net608),
    .X(clknet_1_1__leaf_net608));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net600 (.A(net600),
    .X(clknet_0_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net600 (.A(clknet_0_net600),
    .X(clknet_1_0__leaf_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net600 (.A(clknet_0_net600),
    .X(clknet_1_1__leaf_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net711 (.A(net711),
    .X(clknet_0_net711));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net711 (.A(clknet_0_net711),
    .X(clknet_1_0__leaf_net711));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net711 (.A(clknet_0_net711),
    .X(clknet_1_1__leaf_net711));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net611 (.A(net611),
    .X(clknet_0_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net611 (.A(clknet_0_net611),
    .X(clknet_1_0__leaf_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net611 (.A(clknet_0_net611),
    .X(clknet_1_1__leaf_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net577 (.A(net577),
    .X(clknet_0_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net577 (.A(clknet_0_net577),
    .X(clknet_1_0__leaf_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net577 (.A(clknet_0_net577),
    .X(clknet_1_1__leaf_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net798 (.A(net798),
    .X(clknet_0_net798));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net798 (.A(clknet_0_net798),
    .X(clknet_1_0__leaf_net798));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net798 (.A(clknet_0_net798),
    .X(clknet_1_1__leaf_net798));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net511 (.A(net511),
    .X(clknet_0_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net511 (.A(clknet_0_net511),
    .X(clknet_1_0__leaf_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net511 (.A(clknet_0_net511),
    .X(clknet_1_1__leaf_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net797 (.A(net797),
    .X(clknet_0_net797));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net797 (.A(clknet_0_net797),
    .X(clknet_1_0__leaf_net797));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net797 (.A(clknet_0_net797),
    .X(clknet_1_1__leaf_net797));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net602 (.A(net602),
    .X(clknet_0_net602));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net602 (.A(clknet_0_net602),
    .X(clknet_1_0__leaf_net602));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net602 (.A(clknet_0_net602),
    .X(clknet_1_1__leaf_net602));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net495 (.A(net495),
    .X(clknet_0_net495));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net495 (.A(clknet_0_net495),
    .X(clknet_1_0__leaf_net495));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net495 (.A(clknet_0_net495),
    .X(clknet_1_1__leaf_net495));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net502 (.A(net502),
    .X(clknet_0_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net502 (.A(clknet_0_net502),
    .X(clknet_1_0__leaf_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net502 (.A(clknet_0_net502),
    .X(clknet_1_1__leaf_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net796 (.A(net796),
    .X(clknet_0_net796));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net796 (.A(clknet_0_net796),
    .X(clknet_1_0__leaf_net796));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net796 (.A(clknet_0_net796),
    .X(clknet_1_1__leaf_net796));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net777 (.A(net777),
    .X(clknet_0_net777));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net777 (.A(clknet_0_net777),
    .X(clknet_1_0__leaf_net777));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net777 (.A(clknet_0_net777),
    .X(clknet_1_1__leaf_net777));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net398 (.A(net398),
    .X(clknet_0_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_0__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_1__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net610 (.A(net610),
    .X(clknet_0_net610));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net610 (.A(clknet_0_net610),
    .X(clknet_1_0__leaf_net610));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net610 (.A(clknet_0_net610),
    .X(clknet_1_1__leaf_net610));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net420 (.A(net420),
    .X(clknet_0_net420));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net420 (.A(clknet_0_net420),
    .X(clknet_1_0__leaf_net420));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net420 (.A(clknet_0_net420),
    .X(clknet_1_1__leaf_net420));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net391 (.A(net391),
    .X(clknet_0_net391));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net391 (.A(clknet_0_net391),
    .X(clknet_1_0__leaf_net391));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net391 (.A(clknet_0_net391),
    .X(clknet_1_1__leaf_net391));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net389 (.A(net389),
    .X(clknet_0_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_0__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_1__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net776 (.A(net776),
    .X(clknet_0_net776));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net776 (.A(clknet_0_net776),
    .X(clknet_1_0__leaf_net776));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net776 (.A(clknet_0_net776),
    .X(clknet_1_1__leaf_net776));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net775 (.A(net775),
    .X(clknet_0_net775));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net775 (.A(clknet_0_net775),
    .X(clknet_1_0__leaf_net775));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net775 (.A(clknet_0_net775),
    .X(clknet_1_1__leaf_net775));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net595 (.A(net595),
    .X(clknet_0_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_0__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_1__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net901 (.A(net901),
    .X(clknet_0_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net901 (.A(clknet_0_net901),
    .X(clknet_1_0__leaf_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net901 (.A(clknet_0_net901),
    .X(clknet_1_1__leaf_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net186 (.A(net186),
    .X(clknet_0_net186));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net186 (.A(clknet_0_net186),
    .X(clknet_1_0__leaf_net186));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net186 (.A(clknet_0_net186),
    .X(clknet_1_1__leaf_net186));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net910 (.A(net910),
    .X(clknet_0_net910));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net910 (.A(clknet_0_net910),
    .X(clknet_1_0__leaf_net910));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net910 (.A(clknet_0_net910),
    .X(clknet_1_1__leaf_net910));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net179 (.A(net179),
    .X(clknet_0_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_0__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_1__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net180 (.A(net180),
    .X(clknet_0_net180));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net180 (.A(clknet_0_net180),
    .X(clknet_1_0__leaf_net180));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net180 (.A(clknet_0_net180),
    .X(clknet_1_1__leaf_net180));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net759 (.A(net759),
    .X(clknet_0_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net759 (.A(clknet_0_net759),
    .X(clknet_1_0__leaf_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net759 (.A(clknet_0_net759),
    .X(clknet_1_1__leaf_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net924 (.A(net924),
    .X(clknet_0_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net924 (.A(clknet_0_net924),
    .X(clknet_1_0__leaf_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net924 (.A(clknet_0_net924),
    .X(clknet_1_1__leaf_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net905 (.A(net905),
    .X(clknet_0_net905));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net905 (.A(clknet_0_net905),
    .X(clknet_1_0__leaf_net905));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net905 (.A(clknet_0_net905),
    .X(clknet_1_1__leaf_net905));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net177 (.A(net177),
    .X(clknet_0_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net177 (.A(clknet_0_net177),
    .X(clknet_1_0__leaf_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net177 (.A(clknet_0_net177),
    .X(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net902 (.A(net902),
    .X(clknet_0_net902));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net902 (.A(clknet_0_net902),
    .X(clknet_1_0__leaf_net902));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net902 (.A(net1046),
    .X(clknet_1_1__leaf_net902));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net709 (.A(net709),
    .X(clknet_0_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net709 (.A(clknet_0_net709),
    .X(clknet_1_0__leaf_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net709 (.A(clknet_0_net709),
    .X(clknet_1_1__leaf_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net758 (.A(net758),
    .X(clknet_0_net758));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net758 (.A(clknet_0_net758),
    .X(clknet_1_0__leaf_net758));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net758 (.A(clknet_0_net758),
    .X(clknet_1_1__leaf_net758));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net281 (.A(net281),
    .X(clknet_0_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net281 (.A(clknet_0_net281),
    .X(clknet_1_0__leaf_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net281 (.A(clknet_0_net281),
    .X(clknet_1_1__leaf_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net911 (.A(net911),
    .X(clknet_0_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net911 (.A(clknet_0_net911),
    .X(clknet_1_0__leaf_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net911 (.A(clknet_0_net911),
    .X(clknet_1_1__leaf_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net276 (.A(net276),
    .X(clknet_0_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net276 (.A(clknet_0_net276),
    .X(clknet_1_0__leaf_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net276 (.A(clknet_0_net276),
    .X(clknet_1_1__leaf_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net170 (.A(net170),
    .X(clknet_0_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net170 (.A(clknet_0_net170),
    .X(clknet_1_0__leaf_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net170 (.A(clknet_0_net170),
    .X(clknet_1_1__leaf_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net744 (.A(net744),
    .X(clknet_0_net744));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net744 (.A(clknet_0_net744),
    .X(clknet_1_0__leaf_net744));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net744 (.A(clknet_0_net744),
    .X(clknet_1_1__leaf_net744));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net532 (.A(net532),
    .X(clknet_0_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net532 (.A(clknet_0_net532),
    .X(clknet_1_0__leaf_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net532 (.A(clknet_0_net532),
    .X(clknet_1_1__leaf_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net879 (.A(net879),
    .X(clknet_0_net879));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net879 (.A(clknet_0_net879),
    .X(clknet_1_0__leaf_net879));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net879 (.A(clknet_0_net879),
    .X(clknet_1_1__leaf_net879));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net710 (.A(net710),
    .X(clknet_0_net710));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net710 (.A(clknet_0_net710),
    .X(clknet_1_0__leaf_net710));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net710 (.A(clknet_0_net710),
    .X(clknet_1_1__leaf_net710));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net19),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net1025),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net19),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net1027),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net1032),
    .X(net1029));
 sky130_fd_sc_hd__buf_2 rebuffer6 (.A(net884),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net1),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net21),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net1032),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net23),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net155),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net1035),
    .X(net1036));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer13 (.A(net171),
    .X(net1037));
 sky130_fd_sc_hd__clkbuf_1 clone14 (.A(net22),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net22),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net1041),
    .X(net1040));
 sky130_fd_sc_hd__clkbuf_1 clone17 (.A(net922),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net36),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net1042),
    .X(net1043));
 sky130_fd_sc_hd__clkbuf_1 clone20 (.A(net971),
    .X(net1044));
 sky130_fd_sc_hd__clkbuf_1 clone21 (.A(net17),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(clknet_0_net902),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net799),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net816),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net753),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net727),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net757),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net346),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net792),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net453),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net699),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net921),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net764),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net772),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net435),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net805),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net432),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net769),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net809),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net800),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net735),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net747),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net986),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net770),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net676),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net734),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net704),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net698),
    .X(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_C (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A2 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A0 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_B (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_X (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_S0 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_C (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_A (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_A (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_X (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A2 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_B (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_S0 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_B (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_X (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_C1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A3 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_X (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A3 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_X (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A0 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_X (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A3 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_X (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A0 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_SCD (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_C (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_C (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_C (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_X (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A0 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_D1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_C_N (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_X (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_S1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_X (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_S0 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A0 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S0 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_X (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A0 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A3 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S0 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_SCD (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_C1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_X (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_S0 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_X (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A3 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A0 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_C1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_X (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_X (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A0 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_SCD (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_X (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A0 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S0 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_X (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A3 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A3 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_X (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_X (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_S0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_D (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_X (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_C1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_Q_N (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A1 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A1 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S0 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A1 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A2 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_S1 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_B1 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_X (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A0 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_X (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A0 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_S1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A0 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_X (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A3 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A3 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_Q_N (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_X (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S0 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A3 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S0 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_S1 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A3 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_X (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_X (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_C1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A3 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_X (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_C1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_B1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_B1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_X (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A3 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_C1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_C (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_D1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A3 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_X (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_C1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_X (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_D_N (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A0 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_X (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_X (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A0 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A3 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_D1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_S0 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_S0 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_X (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_B (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_B1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_S1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_C (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_X (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A0 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A3 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_X (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A0 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_X (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_X (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_S0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A0 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_X (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A2 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A2 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_C (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_A (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_C1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_B (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A0 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_D1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_X (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_D1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_B (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_X (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A0 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_D_N (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_X (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A3 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A0 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A3 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_C (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_X (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A3 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A0 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_S0 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S0 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_D_N (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_X (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_X (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_X (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A3 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S0 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_X (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A0 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_S0 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_B1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A3 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_C_N (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_D1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_X (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A0 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A0 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_B (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_X (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A0 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_X (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S0 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A0 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A0 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_S1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_D_N (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_X (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A0 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_S1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_B (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_X (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A2 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_S1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_C_N (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_C_N (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_X (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A3 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_C (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_C1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_X (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_C_N (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_X (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_C_N (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_X (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A0 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_X (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A0 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_RESET_B (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A0 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_X (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer10_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A2 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_X (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A0 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A2 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A3 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A3 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A3 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_C_N (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_X (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_S0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_C1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_Q_N (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_Q (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A0 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_X (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A0 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_S0 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_X (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A3 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_X (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A3 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A3 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_X (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A0 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A2 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A2 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A0 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_X (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_C (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_X (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A3 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A3 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_X (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A0 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A3 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_X (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A0 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S0 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A0 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S0 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_X (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A3 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A3 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_X (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S0 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A3 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_X (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A0 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S0 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S0 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_X (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S0 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A0 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S0 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_X (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_X (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_X (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A0 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_SCD (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_C (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_X (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A3 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A3 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_B (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_X (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_X (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A3 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A0 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_B1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_B1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_C (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_X (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_B1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_RESET_B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_X (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S0 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A0 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_X (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A0 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A3 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_X (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A0 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_X (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_X (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A0 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_SET_B (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A0 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_S0 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A2 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A2 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_B (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_X (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A0 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A3 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A0 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_X (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A0 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A3 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A2 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A2 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A3 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_S0 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_X (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A2 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_D (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_X (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_X (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A0 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_D1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_X (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A0 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A2 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_X (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A0 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A3 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_X (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A0 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_B (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_X (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_X (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A3 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_SCE (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_C1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_X (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A2 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A3 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_X (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A0 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_RESET_B (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_SCD (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_RESET_B (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_X (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A2 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A3 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_X (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A3 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A0 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A2 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_S0 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_X (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold28_A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A3 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S0 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S0 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A3 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_Q_N (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A0 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A2 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_B (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_Q (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_X (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A0 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_S0 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A3 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_C_N (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A0 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A3 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A2 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A3 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_X (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer18_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_X (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A0 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A0 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_X (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A2 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A3 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A3 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A0 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_X (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_D (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_X (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_SCD (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_C (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_X (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_X (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A2 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_X (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A1 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A2 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_B1 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_S1 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_C1 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_X (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S1 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A3 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A1 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A1 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_X (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A3 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_C1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_D1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_X (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A0 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_SCD (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_B (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_S0 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_X (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A1 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_S0 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A0 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A3 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A3 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_S0 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_X (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A0 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A3 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_SCE (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_B1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_X (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A0 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_X (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A3 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_X (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A3 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A3 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_SCD (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_B1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_C1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_X (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A0 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_X (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A0 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A2 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S0 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A1 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_RESET_B (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_X (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A0 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S1 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A2 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_X (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A3 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_X (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A0 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A1 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_X (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A0 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_X (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_SCE (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_X (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_X (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A0 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_S0 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_C (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_X (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A0 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_X (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A0 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A2 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_X (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A0 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_Q (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A0 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A2 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_D1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_X (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A0 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A0 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A3 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_SCD (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_X (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A2 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A2 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_X (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A1 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A0 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_X (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A1 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_X (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A2 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A3 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A0 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A3 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A3 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_X (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_D (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_X (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_C (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_X (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_S0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A3 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A3 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_D (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_X (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_Q (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S0 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S0 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_S0 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_S0 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_S0 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_B1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_Q_N (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_SCE (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_S0 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_X (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold45_A (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_Q_N (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S0 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S0 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A3 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_C_N (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_C_N (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_SET_B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_C (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_X (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_Q (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S0 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S0 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A2 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S0 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_C_N (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S0 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_Q (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S1 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_Q (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold48_A (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_Q (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S0 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S0 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S0 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_C1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_C1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_D1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold31_A (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_Q (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S0 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S0 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S0 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_D1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_X (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold47_A (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_Q (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S0 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_S1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_X (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_Q (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A3 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S1 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_S1 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_Q_N (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S1 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S0 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_X (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_S1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_D1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S0 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S0 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge860_Q_N (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A3 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_Q (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A2 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S0 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_X (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold41_A (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_Q (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S0 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A3 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_Q (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S1 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S0 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_Q (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_S1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S0 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_Q (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S1 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S1 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S0 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_S0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_S1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_X (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_Q (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S0 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A3 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge885_Q (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S1 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S0 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_Q (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_S0 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_S0 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_S0 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_Q (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_SET_B (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_D1 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_C1 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_D1 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_Q (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_S0 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_S0 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_X (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_Q (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S0 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S0 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_Q_N (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_S0 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_Q (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_S0 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap172_A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_Q (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S0 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_Q_N (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A3 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S0 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold34_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_Q (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S0 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_S1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S0 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_Q (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_S1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_S1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_C (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_X (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_Q (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_S0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A3 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A3 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_S0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A3 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_D1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_S1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_Q (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_S0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_D1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_X (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_Q (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S0 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_S0 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_s922_Q (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_S1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A3 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_X (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A3 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_S0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_B (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_X (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_Q_N (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_Q (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_S0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_Q (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_Q (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S0 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_S0 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_D1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_C (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A3 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_Q (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S0 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A2 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A3 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_X (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_SCE (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A3 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_C (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_SCE (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_RESET_B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_S0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_X (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_C (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_X (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_SCE (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A3 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_A1 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_B (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_RESET_B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_X (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_D1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_X (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_C1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_C1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_X (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A0 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A0 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A0 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A3 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_D1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_X (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A0 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_B (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A2 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A3 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A0 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_A (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A3 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A3 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A1 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_S0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A3 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A2 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_A (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A2 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A2 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_B (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A3 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A3 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A2 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A3 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_A (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A3 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A2 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_D1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_A (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A3 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_S1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_B1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_C1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_C1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_S1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_C_N (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A3 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A2 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_B1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A2 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_D_N (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_C1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A3 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_A (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_C1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_B (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_C (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_B1 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A2 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A2 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_C1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_S0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_C1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_B1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_A (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A0 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A3 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_C1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_X (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A3 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A2 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_C1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_S0 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A3 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_D (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_C (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_D1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_C1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A3 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_S0 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A2 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_B1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_C_N (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_D1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_C (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A2 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_C (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A2 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A0 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A2 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_C1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A1 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_B (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_D_N (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A2 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_D_N (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_X (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_B (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_B (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A2 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A0 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_D1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_C (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_B (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A2 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_B1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_B (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_S1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S0 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A3 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A0 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_S0 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_C (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A2 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S0 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A2 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S0 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A0 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A0 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A2 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A3 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A2 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_B (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A3 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A3 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_B (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_A (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A3 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A3 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A2 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_B1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_D1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_C_N (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_D_N (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_X (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_B (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_C (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_C (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_B (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_B1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S1 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A0 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_S0 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_B (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_X (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A0 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A3 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A1 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A0 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A1 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_B (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A0 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A2 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_X (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_B (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A3 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A0 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A1 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A2 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_C1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_X (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_RESET_B (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_C (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A1 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A3 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_X (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A3 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_Q (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A3 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_S0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_A3 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_A1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A3 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A3 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A3 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_D1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_X (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_X (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S0 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_RESET_B (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_X (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A3 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S0 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A3 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A3 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_X (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A1 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer6_A (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A3 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A2 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A2 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_X (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A2 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A3 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_Q (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_S0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A2 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A2 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_SCE (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_B (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_B (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_X (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A2 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_X (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A0 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A2 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A2 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A2 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_X (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_Q (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A3 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_S0 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A2 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_X (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge875_Q (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A3 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_S0 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_Q (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_Q_N (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_S0 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_S0 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A3 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_S0 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A2 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A2 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_Q (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_Q (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_S0 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_D1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_S0 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A2 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A3 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_X (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_Q (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S0 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_X (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A2 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A2 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A2 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_Q (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge832_Q (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A1 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A3 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_X (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_D (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_X (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_X (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S1 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A3 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_Q (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A1 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A2 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_X (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A2 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A2 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_X (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A3 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_S0 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_X (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold32_A (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_Q (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A3 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A2 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_X (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_Q (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_S1 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S0 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A3 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A2 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_C_N (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_X (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_X (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_SCE (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_B1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_C_N (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A3 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_SET_B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A2 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_C (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_X (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_X (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_RESET_B (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_S0 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A2 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A0 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A3 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_X (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A2 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_B1 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_S0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A2 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_X (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A2 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A2 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_D_N (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_X (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_SCE (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_C1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A3 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A3 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_C1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_X (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_C1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_C (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_B1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S0 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_X (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_B1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_C_N (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_S1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A3 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A3 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_X (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A0 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A3 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_A1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_SCE (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_C_N (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_B (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_C1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A0 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A2 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_X (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_S1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A3 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A3 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_X (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_SET_B (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_C1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_D_N (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_S1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_X (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A2 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A2 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_S0 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_X (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_B1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A3 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A2 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_C (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A3 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_D1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A3 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A2 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_X (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A0 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_S1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S0 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S0 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_SET_B (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A2 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_D1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A3 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_D_N (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_SCE (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_X (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A0 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_D_N (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A0 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_B (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_B1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_SCD (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_X (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A3 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_B (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A2 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_C_N (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A2 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S0 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_C1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_X (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A0 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A2 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A3 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_C1 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_D_N (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_C (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A3 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A2 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S0 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A0 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_X (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A3 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_S1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A3 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_D1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A3 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_D1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_C (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_X (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_A2 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A2 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_S0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_B1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_S1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A2 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_C1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_C (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_D1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_B1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_X (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A2 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A3 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_S0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_S0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A3 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_X (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_C (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_S1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_S1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_SCD (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_S0 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_B1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A3 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_S0 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_X (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_C1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S0 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_S0 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S0 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_X (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_S0 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A0 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A3 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_X (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_C_N (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_S0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_B1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_D1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_X (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_S0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A3 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_C1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_X (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_C1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_C_N (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_C_N (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_X (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_C (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_D1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_C (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_B1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_B1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_S1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_C (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_X (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_B (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_C1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_D_N (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_S0 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_D1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S0 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_X (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_SCE (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_D (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_D_N (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_D1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_D_N (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_C_N (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_S0 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_D_N (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_C (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_X (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_S1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A0 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A3 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_X (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_B1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_S1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S0 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_C1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_C (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_C1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_X (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_S0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_C1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A3 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_B1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A3 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_C1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_B (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_X (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A2 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S0 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_B1 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_RESET_B (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_C1 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_B1 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A1 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_C1 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_B (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone20_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_X (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_S0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_C1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_S0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_X (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_S0 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_S0 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_C (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_S1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_B1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_C (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A3 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_D_N (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A2 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_X (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_S0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_D1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_C (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A2 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_B (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_B (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_X (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A3 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_S0 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A3 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A0 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A3 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A2 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_X (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_C (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A3 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A2 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A3 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_C_N (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_A2 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_C_N (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_C1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_X (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S0 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A3 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_S0 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_A (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_X (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_C (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_S0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_C (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_C (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_C1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_C (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_D1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A2 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_X (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_S0 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_SCE (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_D1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_S1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_D1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_D1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_S0 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_D_N (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_X (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A3 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A2 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_X (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_S0 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_S0 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A2 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_C1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_S1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A0 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_X (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_S1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_C (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_S0 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_C (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_C (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A0 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_X (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_S0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold43_A (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_X (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_S1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A3 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_D1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_S1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_S1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_D1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_D1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap172_X (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_X (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_S0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A3 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_B1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_D1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A3 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_X (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_C1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A3 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A3 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_X (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A3 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_C1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_X (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_B1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A3 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A0 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_D1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_C (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_C (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_S0 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_C (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_X (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_C (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_S1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A2 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A3 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A2 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A3 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_X (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S0 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_X (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A3 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A3 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_C (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_X (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_C_N (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_D1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_D1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A2 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_C (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_C (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_X (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_C1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_D1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_B1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A3 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A0 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_X (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_S0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_S0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A3 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A3 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A3 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_X (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_D1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_S1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_D_N (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_S0 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_C (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_S0 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_D1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_C (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_X (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_D1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_S1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_D_N (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_S1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_C1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_D_N (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_X (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A3 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A3 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_S0 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_SCE (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_D1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_C (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_X (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S0 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_C_N (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_C_N (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_X (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A3 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_C1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A3 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A2 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S0 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A2 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_C1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_X (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_C_N (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A0 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_C (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_D1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_C (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_X (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_D1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_S0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_X (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S0 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_S0 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_S1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A0 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A3 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_S0 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_B (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_X (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_D1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_C (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A3 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_S1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_C1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_D_N (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_X (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_D_N (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A3 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_C1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_RESET_B (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_C (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_D1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_X (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_C1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A3 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_B (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A3 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_SCD (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_X (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A2 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_C1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_C1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_C (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_B1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_C_N (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_X (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_A (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_B (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A2 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_S0 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_X (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A2 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A0 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_S1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_C (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_X (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_C1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_S0 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_C_N (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_C1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_D_N (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_X (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_C (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_S1 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_C (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_C (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A2 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_X (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A3 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_C1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_D1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_S0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_B1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_X (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_C (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_D1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_X (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_S0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_X (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_S0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_C1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_C (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_S1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A3 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A3 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_X (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A2 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_C_N (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_C_N (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_C1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_X (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A0 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_X (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_A2 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A2 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_S0 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_C (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_S0 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_X (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_D_N (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_D1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_B1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_D1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A2 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_C1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_D1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_C (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_X (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_S0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_D1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_B (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_X (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A3 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_S0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A3 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_S0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_B (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_X (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_D_N (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_B (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A3 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A2 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A2 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_SLEEP_B (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s929_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge885_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s921_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s933_SLEEP_B (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s935_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_GATE (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_GATE (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_SLEEP_B (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s905_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s922_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s924_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s938_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s939_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s940_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_GATE (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge875_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s908_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge877_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s926_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge864_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge848_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s910_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_GATE (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge847_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_GATE (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_GATE (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_X (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S1 (.DIODE(clknet_1_1__leaf_net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S1 (.DIODE(clknet_1_1__leaf_net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(clknet_1_1__leaf_net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net775_X (.DIODE(clknet_1_1__leaf_net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_S1 (.DIODE(clknet_1_1__leaf_net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_S1 (.DIODE(clknet_1_1__leaf_net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_S1 (.DIODE(clknet_1_1__leaf_net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(clknet_1_1__leaf_net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net901_X (.DIODE(clknet_1_1__leaf_net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_A (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_X (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer6_X (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer16_A (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_SCE (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_S1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S0 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone17_X (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_C1 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A3 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_S1 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A3 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone21_X (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net1011));
 sky130_fd_sc_hd__mux4_1 clone1 (.A0(net842),
    .A1(net112),
    .A2(net123),
    .A3(net1009),
    .S0(net971),
    .S1(net957),
    .X(net1073));
 sky130_fd_sc_hd__and3_1 clone2 (.A(net1),
    .B(net860),
    .C(net0),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net82),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net1075),
    .X(net1076));
 sky130_fd_sc_hd__mux4_1 clone18 (.A0(net862),
    .A1(net860),
    .A2(net840),
    .A3(net871),
    .S0(net990),
    .S1(net858),
    .X(net1077));
 sky130_fd_sc_hd__mux4_1 clone19 (.A0(net102),
    .A1(net100),
    .A2(net827),
    .A3(net104),
    .S0(net97),
    .S1(net949),
    .X(net1078));
 sky130_fd_sc_hd__mux4_1 clone22 (.A0(net842),
    .A1(net112),
    .A2(net123),
    .A3(net1009),
    .S0(net971),
    .S1(net957),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net880),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net880),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net1081),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net1081),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(net1083),
    .X(net1084));
 sky130_fd_sc_hd__a2111o_1 clone28 (.A1(net951),
    .A2(net884),
    .B1(net664),
    .C1(net754),
    .D1(net755),
    .X(net1085));
 sky130_fd_sc_hd__a2111o_1 clone29 (.A1(net16),
    .A2(net18),
    .B1(net970),
    .C1(net13),
    .D1(net19),
    .X(net1086));
 sky130_fd_sc_hd__or4bb_1 clone30 (.A(net8),
    .B(net6),
    .C_N(net970),
    .D_N(net951),
    .X(net1087));
 sky130_fd_sc_hd__buf_2 rebuffer31 (.A(net98),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(net1088),
    .X(net1089));
 sky130_fd_sc_hd__a2111o_1 clone33 (.A1(net28),
    .A2(net871),
    .B1(net42),
    .C1(net856),
    .D1(net43),
    .X(net1090));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
