module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in62,
    in63,
    in64,
    in65,
    in66,
    in67,
    in68,
    in69,
    in7,
    in70,
    in71,
    in72,
    in73,
    in74,
    in75,
    in76,
    in77,
    in78,
    in79,
    in8,
    in80,
    in81,
    in82,
    in83,
    in84,
    in85,
    in86,
    in87,
    in88,
    in89,
    in9,
    in90,
    in91,
    in92,
    in93,
    in94,
    in95,
    in96,
    in97,
    in98,
    in99,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out62,
    out63,
    out64,
    out65,
    out66,
    out67,
    out68,
    out69,
    out7,
    out70,
    out71,
    out72,
    out73,
    out74,
    out75,
    out76,
    out77,
    out78,
    out79,
    out8,
    out80,
    out81,
    out82,
    out83,
    out84,
    out85,
    out86,
    out87,
    out88,
    out89,
    out9,
    out90,
    out91,
    out92,
    out93,
    out94,
    out95,
    out96,
    out97,
    out98,
    out99,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in62;
 input in63;
 input in64;
 input in65;
 input in66;
 input in67;
 input in68;
 input in69;
 input in7;
 input in70;
 input in71;
 input in72;
 input in73;
 input in74;
 input in75;
 input in76;
 input in77;
 input in78;
 input in79;
 input in8;
 input in80;
 input in81;
 input in82;
 input in83;
 input in84;
 input in85;
 input in86;
 input in87;
 input in88;
 input in89;
 input in9;
 input in90;
 input in91;
 input in92;
 input in93;
 input in94;
 input in95;
 input in96;
 input in97;
 input in98;
 input in99;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out62;
 output out63;
 output out64;
 output out65;
 output out66;
 output out67;
 output out68;
 output out69;
 output out7;
 output out70;
 output out71;
 output out72;
 output out73;
 output out74;
 output out75;
 output out76;
 output out77;
 output out78;
 output out79;
 output out8;
 output out80;
 output out81;
 output out82;
 output out83;
 output out84;
 output out85;
 output out86;
 output out87;
 output out88;
 output out89;
 output out9;
 output out90;
 output out91;
 output out92;
 output out93;
 output out94;
 output out95;
 output out96;
 output out97;
 output out98;
 output out99;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net182;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_0_net615;
 wire clknet_1_0__leaf_net615;
 wire clknet_1_1__leaf_net615;
 wire clknet_0_net475;
 wire clknet_1_0__leaf_net475;
 wire clknet_1_1__leaf_net475;
 wire clknet_0_net799;
 wire clknet_1_0__leaf_net799;
 wire clknet_1_1__leaf_net799;
 wire clknet_0_net370;
 wire clknet_1_0__leaf_net370;
 wire clknet_1_1__leaf_net370;
 wire clknet_0_net512;
 wire clknet_1_0__leaf_net512;
 wire clknet_1_1__leaf_net512;
 wire clknet_0_net295;
 wire clknet_1_0__leaf_net295;
 wire clknet_1_1__leaf_net295;
 wire clknet_0_net400;
 wire clknet_1_0__leaf_net400;
 wire clknet_1_1__leaf_net400;
 wire clknet_0_net300;
 wire clknet_1_0__leaf_net300;
 wire clknet_1_1__leaf_net300;
 wire clknet_0_net289;
 wire clknet_1_0__leaf_net289;
 wire clknet_1_1__leaf_net289;
 wire clknet_0_net305;
 wire clknet_1_0__leaf_net305;
 wire clknet_1_1__leaf_net305;
 wire clknet_0_net301;
 wire clknet_1_0__leaf_net301;
 wire clknet_1_1__leaf_net301;
 wire clknet_0_net268;
 wire clknet_1_0__leaf_net268;
 wire clknet_1_1__leaf_net268;
 wire clknet_0_net255;
 wire clknet_1_0__leaf_net255;
 wire clknet_1_1__leaf_net255;
 wire clknet_0_net614;
 wire clknet_1_0__leaf_net614;
 wire clknet_1_1__leaf_net614;
 wire clknet_0_net473;
 wire clknet_1_0__leaf_net473;
 wire clknet_1_1__leaf_net473;
 wire clknet_0_net793;
 wire clknet_1_0__leaf_net793;
 wire clknet_1_1__leaf_net793;
 wire clknet_0_net367;
 wire clknet_1_0__leaf_net367;
 wire clknet_1_1__leaf_net367;
 wire clknet_0_net198;
 wire clknet_1_0__leaf_net198;
 wire clknet_1_1__leaf_net198;
 wire clknet_0_net199;
 wire clknet_1_0__leaf_net199;
 wire clknet_1_1__leaf_net199;
 wire clknet_0_net200;
 wire clknet_1_0__leaf_net200;
 wire clknet_1_1__leaf_net200;
 wire clknet_0_net179;
 wire clknet_1_0__leaf_net179;
 wire clknet_1_1__leaf_net179;
 wire clknet_0_net178;
 wire clknet_1_0__leaf_net178;
 wire clknet_1_1__leaf_net178;
 wire clknet_0_net375;
 wire clknet_1_0__leaf_net375;
 wire clknet_1_1__leaf_net375;
 wire clknet_0_net277;
 wire clknet_1_0__leaf_net277;
 wire clknet_1_1__leaf_net277;
 wire clknet_0_net281;
 wire clknet_1_0__leaf_net281;
 wire clknet_1_1__leaf_net281;
 wire clknet_0_net282;
 wire clknet_1_0__leaf_net282;
 wire clknet_1_1__leaf_net282;
 wire clknet_0_net276;
 wire clknet_1_0__leaf_net276;
 wire clknet_1_1__leaf_net276;
 wire clknet_0_net166;
 wire clknet_1_0__leaf_net166;
 wire clknet_1_1__leaf_net166;
 wire clknet_0_net769;
 wire clknet_1_0__leaf_net769;
 wire clknet_1_1__leaf_net769;
 wire clknet_0_net162;
 wire clknet_1_0__leaf_net162;
 wire clknet_1_1__leaf_net162;
 wire clknet_0_net161;
 wire clknet_1_0__leaf_net161;
 wire clknet_1_1__leaf_net161;
 wire clknet_0_net159;
 wire clknet_1_0__leaf_net159;
 wire clknet_1_1__leaf_net159;
 wire clknet_0_net766;
 wire clknet_1_0__leaf_net766;
 wire clknet_1_1__leaf_net766;
 wire clknet_0_net786;
 wire clknet_1_0__leaf_net786;
 wire clknet_1_1__leaf_net786;
 wire clknet_0_net742;
 wire clknet_1_0__leaf_net742;
 wire clknet_1_1__leaf_net742;
 wire clknet_0_net97;
 wire clknet_1_0__leaf_net97;
 wire clknet_1_1__leaf_net97;
 wire clknet_0_net800;
 wire clknet_1_0__leaf_net800;
 wire clknet_1_1__leaf_net800;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;

 sky130_fd_sc_hd__a21bo_1 c100 (.A1(net695),
    .A2(net715),
    .B1_N(net717),
    .X(net0));
 sky130_fd_sc_hd__a21bo_1 c101 (.A1(net714),
    .A2(net702),
    .B1_N(net663),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c102 (.A0(net632),
    .A1(net673),
    .A2(net720),
    .A3(net700),
    .S0(net703),
    .S1(net716),
    .X(net2));
 sky130_fd_sc_hd__a31o_1 c103 (.A1(net720),
    .A2(net1),
    .A3(net647),
    .B1(net722),
    .X(net774));
 sky130_fd_sc_hd__a21bo_1 c104 (.A1(net711),
    .A2(net662),
    .B1_N(net670),
    .X(net3));
 sky130_fd_sc_hd__a31o_2 c105 (.A1(net713),
    .A2(net649),
    .A3(net719),
    .B1(net3),
    .X(net758));
 sky130_fd_sc_hd__a21bo_1 c106 (.A1(net717),
    .A2(net721),
    .B1_N(net848),
    .X(net4));
 sky130_fd_sc_hd__a41o_1 c107 (.A1(net716),
    .A2(net3),
    .A3(net691),
    .A4(net695),
    .B1(net676),
    .X(net5));
 sky130_fd_sc_hd__a41o_1 c108 (.A1(net2),
    .A2(net720),
    .A3(net716),
    .A4(net758),
    .B1(net712),
    .X(net756));
 sky130_fd_sc_hd__mux4_1 c109 (.A0(net1),
    .A1(net756),
    .A2(net5),
    .A3(net710),
    .S0(net711),
    .S1(net719),
    .X(net6));
 sky130_fd_sc_hd__xnor2_1 c110 (.A(net889),
    .B(net628),
    .Y(net7));
 sky130_fd_sc_hd__xnor2_1 c111 (.A(net636),
    .B(net629),
    .Y(net789));
 sky130_fd_sc_hd__xnor2_2 c112 (.A(net703),
    .B(net704),
    .Y(net791));
 sky130_fd_sc_hd__xnor2_1 c113 (.A(net647),
    .B(net840),
    .Y(net784));
 sky130_fd_sc_hd__xnor2_1 c114 (.A(net719),
    .B(net840),
    .Y(net792));
 sky130_fd_sc_hd__xnor2_1 c115 (.A(net646),
    .B(net0),
    .Y(net8));
 sky130_fd_sc_hd__xnor2_1 c116 (.A(net675),
    .B(net714),
    .Y(net9));
 sky130_fd_sc_hd__a21bo_2 c117 (.A1(net676),
    .A2(net684),
    .B1_N(net636),
    .X(net10));
 sky130_fd_sc_hd__a21bo_1 c118 (.A1(net2),
    .A2(net680),
    .B1_N(net840),
    .X(net798));
 sky130_fd_sc_hd__a21bo_1 c119 (.A1(net8),
    .A2(net6),
    .B1_N(net840),
    .X(net788));
 sky130_fd_sc_hd__a41o_1 c120 (.A1(net10),
    .A2(net718),
    .A3(net632),
    .A4(net712),
    .B1(net798),
    .X(net11));
 sky130_fd_sc_hd__mux4_1 c121 (.A0(net11),
    .A1(net699),
    .A2(net789),
    .A3(net840),
    .S0(net704),
    .S1(net10),
    .X(net12));
 sky130_fd_sc_hd__a21bo_2 c122 (.A1(net638),
    .A2(net704),
    .B1_N(net0),
    .X(net13));
 sky130_fd_sc_hd__a21bo_1 c123 (.A1(net13),
    .A2(net840),
    .B1_N(net10),
    .X(net794));
 sky130_fd_sc_hd__a21bo_1 c124 (.A1(net12),
    .A2(net712),
    .B1_N(net840),
    .X(net802));
 sky130_fd_sc_hd__a41o_1 c125 (.A1(net10),
    .A2(net802),
    .A3(net840),
    .A4(net13),
    .B1(net756),
    .X(net768));
 sky130_fd_sc_hd__a21bo_1 c126 (.A1(net712),
    .A2(net13),
    .B1_N(net718),
    .X(net781));
 sky130_fd_sc_hd__mux4_1 c127 (.A0(net663),
    .A1(net13),
    .A2(net10),
    .A3(net788),
    .S0(net8),
    .S1(net791),
    .X(net775));
 sky130_fd_sc_hd__a21bo_1 c128 (.A1(net0),
    .A2(net781),
    .B1_N(net7),
    .X(net795));
 sky130_fd_sc_hd__a21bo_1 c129 (.A1(net631),
    .A2(net840),
    .B1_N(net775),
    .X(net772));
 sky130_fd_sc_hd__a41o_1 c130 (.A1(net632),
    .A2(net647),
    .A3(net9),
    .A4(net756),
    .B1(net768),
    .X(net14));
 sky130_fd_sc_hd__a21bo_1 c131 (.A1(net718),
    .A2(net10),
    .B1_N(net14),
    .X(net15));
 sky130_fd_sc_hd__xnor2_4 c132 (.A(net657),
    .B(net679),
    .Y(net16));
 sky130_fd_sc_hd__xnor2_4 c133 (.A(net633),
    .B(net852),
    .Y(net17));
 sky130_fd_sc_hd__a21bo_4 c134 (.A1(net851),
    .A2(net633),
    .B1_N(net838),
    .X(net777));
 sky130_fd_sc_hd__a21bo_4 c135 (.A1(net777),
    .A2(net632),
    .B1_N(net849),
    .X(net761));
 sky130_fd_sc_hd__xnor2_4 c136 (.A(net646),
    .B(net17),
    .Y(net18));
 sky130_fd_sc_hd__a21bo_2 c137 (.A1(net646),
    .A2(net633),
    .B1_N(net837),
    .X(net19));
 sky130_fd_sc_hd__xnor2_2 c138 (.A(net17),
    .B(net18),
    .Y(net730));
 sky130_fd_sc_hd__a21bo_4 c139 (.A1(net761),
    .A2(net18),
    .B1_N(net825),
    .X(net20));
 sky130_fd_sc_hd__xnor2_4 c140 (.A(net635),
    .B(net836),
    .Y(net21));
 sky130_fd_sc_hd__a21bo_4 c141 (.A1(net837),
    .A2(net18),
    .B1_N(net632),
    .X(net760));
 sky130_fd_sc_hd__xnor2_2 c142 (.A(net635),
    .B(net636),
    .Y(net22));
 sky130_fd_sc_hd__a21bo_4 c143 (.A1(net847),
    .A2(net21),
    .B1_N(net838),
    .X(net23));
 sky130_fd_sc_hd__mux4_2 c144 (.A0(net777),
    .A1(net630),
    .A2(net760),
    .A3(net18),
    .S0(net23),
    .S1(net837),
    .X(net24));
 sky130_fd_sc_hd__mux4_2 c145 (.A0(net760),
    .A1(net19),
    .A2(net690),
    .A3(net712),
    .S0(net825),
    .S1(net837),
    .X(net744));
 sky130_fd_sc_hd__a21bo_4 c146 (.A1(net760),
    .A2(net630),
    .B1_N(net849),
    .X(net25));
 sky130_fd_sc_hd__mux4_2 c147 (.A0(net24),
    .A1(net20),
    .A2(net23),
    .A3(net760),
    .S0(net19),
    .S1(net837),
    .X(net26));
 sky130_fd_sc_hd__a31o_4 c148 (.A1(net18),
    .A2(net24),
    .A3(net19),
    .B1(net837),
    .X(net783));
 sky130_fd_sc_hd__xnor2_2 c149 (.A(net25),
    .B(net17),
    .Y(net27));
 sky130_fd_sc_hd__mux4_2 c150 (.A0(net20),
    .A1(net820),
    .A2(net712),
    .A3(net633),
    .S0(net825),
    .S1(net837),
    .X(net771));
 sky130_fd_sc_hd__mux4_2 c151 (.A0(net26),
    .A1(net23),
    .A2(net25),
    .A3(net22),
    .S0(net839),
    .S1(net826),
    .X(net740));
 sky130_fd_sc_hd__a41o_4 c152 (.A1(net823),
    .A2(net20),
    .A3(net771),
    .A4(net838),
    .B1(net825),
    .X(net28));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net21),
    .A1(net28),
    .A2(net818),
    .A3(net823),
    .S0(net25),
    .S1(net771),
    .X(net29));
 sky130_fd_sc_hd__a31o_2 c154 (.A1(net655),
    .A2(net642),
    .A3(net651),
    .B1(net644),
    .X(net30));
 sky130_fd_sc_hd__a21bo_1 c155 (.A1(net652),
    .A2(net646),
    .B1_N(net852),
    .X(net31));
 sky130_fd_sc_hd__a21bo_4 c156 (.A1(net637),
    .A2(net712),
    .B1_N(net653),
    .X(net731));
 sky130_fd_sc_hd__a21bo_1 c157 (.A1(net731),
    .A2(net648),
    .B1_N(net831),
    .X(net32));
 sky130_fd_sc_hd__a31o_2 c158 (.A1(net633),
    .A2(net630),
    .A3(net831),
    .B1(net837),
    .X(net33));
 sky130_fd_sc_hd__a41o_2 c159 (.A1(net32),
    .A2(net831),
    .A3(net637),
    .A4(net24),
    .B1(net826),
    .X(net797));
 sky130_fd_sc_hd__a41o_1 c160 (.A1(net24),
    .A2(net634),
    .A3(net731),
    .A4(net837),
    .B1(net831),
    .X(net34));
 sky130_fd_sc_hd__a21bo_4 c161 (.A1(net771),
    .A2(net650),
    .B1_N(net652),
    .X(net35));
 sky130_fd_sc_hd__a41o_2 c162 (.A1(net644),
    .A2(net661),
    .A3(net830),
    .A4(net650),
    .B1(net690),
    .X(net36));
 sky130_fd_sc_hd__a31o_2 c163 (.A1(net797),
    .A2(net34),
    .A3(net32),
    .B1(net826),
    .X(net725));
 sky130_fd_sc_hd__a21bo_2 c164 (.A1(net660),
    .A2(net36),
    .B1_N(net652),
    .X(net37));
 sky130_fd_sc_hd__mux4_2 c165 (.A0(net18),
    .A1(net37),
    .A2(net647),
    .A3(net731),
    .S0(net832),
    .S1(net837),
    .X(net38));
 sky130_fd_sc_hd__mux4_2 c166 (.A0(net630),
    .A1(net30),
    .A2(net654),
    .A3(net644),
    .S0(net35),
    .S1(net831),
    .X(net732));
 sky130_fd_sc_hd__a21bo_2 c167 (.A1(net634),
    .A2(net731),
    .B1_N(net32),
    .X(net780));
 sky130_fd_sc_hd__a41o_4 c168 (.A1(net38),
    .A2(net34),
    .A3(net831),
    .A4(net797),
    .B1(net813),
    .X(net39));
 sky130_fd_sc_hd__a21bo_2 c169 (.A1(net36),
    .A2(net33),
    .B1_N(net813),
    .X(net40));
 sky130_fd_sc_hd__a41o_2 c170 (.A1(net35),
    .A2(net633),
    .A3(net813),
    .A4(net33),
    .B1(net831),
    .X(net41));
 sky130_fd_sc_hd__a21bo_2 c171 (.A1(net40),
    .A2(net712),
    .B1_N(net41),
    .X(net42));
 sky130_fd_sc_hd__a21bo_4 c172 (.A1(net39),
    .A2(net642),
    .B1_N(net826),
    .X(net43));
 sky130_fd_sc_hd__mux4_2 c173 (.A0(net832),
    .A1(net35),
    .A2(net813),
    .A3(net36),
    .S0(net26),
    .S1(net648),
    .X(net44));
 sky130_fd_sc_hd__a41o_4 c174 (.A1(net813),
    .A2(net26),
    .A3(net43),
    .A4(net832),
    .B1(net826),
    .X(net45));
 sky130_fd_sc_hd__mux4_2 c175 (.A0(net44),
    .A1(net45),
    .A2(net41),
    .A3(net43),
    .S0(net651),
    .S1(net639),
    .X(net803));
 sky130_fd_sc_hd__mux4_2 c176 (.A0(net648),
    .A1(net678),
    .A2(net813),
    .A3(net654),
    .S0(net653),
    .S1(net803),
    .X(net46));
 sky130_fd_sc_hd__a21bo_4 c177 (.A1(net643),
    .A2(net683),
    .B1_N(net761),
    .X(net47));
 sky130_fd_sc_hd__a21bo_1 c178 (.A1(net648),
    .A2(net47),
    .B1_N(net831),
    .X(net48));
 sky130_fd_sc_hd__a21bo_2 c179 (.A1(net24),
    .A2(net38),
    .B1_N(net630),
    .X(net49));
 sky130_fd_sc_hd__a21bo_2 c180 (.A1(net630),
    .A2(net671),
    .B1_N(net47),
    .X(net796));
 sky130_fd_sc_hd__a21bo_1 c181 (.A1(net639),
    .A2(net658),
    .B1_N(net24),
    .X(net50));
 sky130_fd_sc_hd__a21bo_2 c182 (.A1(net30),
    .A2(net50),
    .B1_N(net34),
    .X(net51));
 sky130_fd_sc_hd__a21bo_1 c183 (.A1(net760),
    .A2(net666),
    .B1_N(net643),
    .X(net52));
 sky130_fd_sc_hd__mux4_2 c184 (.A0(net669),
    .A1(net50),
    .A2(net52),
    .A3(net667),
    .S0(net43),
    .S1(net46),
    .X(net53));
 sky130_fd_sc_hd__mux4_2 c185 (.A0(net656),
    .A1(net678),
    .A2(net51),
    .A3(net30),
    .S0(net38),
    .S1(net666),
    .X(net54));
 sky130_fd_sc_hd__a31o_1 c186 (.A1(net49),
    .A2(net680),
    .A3(net682),
    .B1(net54),
    .X(net55));
 sky130_fd_sc_hd__a21bo_4 c187 (.A1(net796),
    .A2(net53),
    .B1_N(net833),
    .X(net728));
 sky130_fd_sc_hd__a21bo_2 c188 (.A1(net646),
    .A2(net649),
    .B1_N(net833),
    .X(net56));
 sky130_fd_sc_hd__mux4_2 c189 (.A0(net41),
    .A1(net56),
    .A2(net728),
    .A3(net669),
    .S0(net683),
    .S1(net639),
    .X(net57));
 sky130_fd_sc_hd__a21bo_1 c190 (.A1(net864),
    .A2(net682),
    .B1_N(net674),
    .X(net58));
 sky130_fd_sc_hd__mux4_2 c191 (.A0(net632),
    .A1(net728),
    .A2(net58),
    .A3(net662),
    .S0(net52),
    .S1(net832),
    .X(net782));
 sky130_fd_sc_hd__a21bo_2 c192 (.A1(net27),
    .A2(net55),
    .B1_N(net832),
    .X(net59));
 sky130_fd_sc_hd__mux4_2 c193 (.A0(net782),
    .A1(net796),
    .A2(net659),
    .A3(net653),
    .S0(net55),
    .S1(net662),
    .X(net60));
 sky130_fd_sc_hd__a41o_2 c194 (.A1(net52),
    .A2(net58),
    .A3(net60),
    .A4(net59),
    .B1(net832),
    .X(net61));
 sky130_fd_sc_hd__a31o_1 c195 (.A1(net54),
    .A2(net58),
    .A3(net850),
    .B1(net59),
    .X(net62));
 sky130_fd_sc_hd__mux4_2 c196 (.A0(net59),
    .A1(net648),
    .A2(net62),
    .A3(net796),
    .S0(net728),
    .S1(net58),
    .X(net63));
 sky130_fd_sc_hd__mux4_2 c197 (.A0(net46),
    .A1(net62),
    .A2(net60),
    .A3(net58),
    .S0(net54),
    .S1(net832),
    .X(net64));
 sky130_fd_sc_hd__a21bo_2 c198 (.A1(net35),
    .A2(net26),
    .B1_N(net638),
    .X(net65));
 sky130_fd_sc_hd__a21bo_4 c199 (.A1(net50),
    .A2(net761),
    .B1_N(net831),
    .X(net66));
 sky130_fd_sc_hd__a41o_1 c200 (.A1(net712),
    .A2(net697),
    .A3(net685),
    .A4(net839),
    .B1(net834),
    .X(net67));
 sky130_fd_sc_hd__a21bo_4 c201 (.A1(net689),
    .A2(net803),
    .B1_N(net777),
    .X(net68));
 sky130_fd_sc_hd__a21bo_1 c202 (.A1(net65),
    .A2(net691),
    .B1_N(net704),
    .X(net69));
 sky130_fd_sc_hd__a21bo_1 c203 (.A1(net66),
    .A2(net698),
    .B1_N(net47),
    .X(net70));
 sky130_fd_sc_hd__mux4_2 c204 (.A0(net678),
    .A1(net45),
    .A2(net66),
    .A3(net797),
    .S0(net850),
    .S1(net810),
    .X(net71));
 sky130_fd_sc_hd__a21bo_4 c205 (.A1(net71),
    .A2(net60),
    .B1_N(net680),
    .X(net746));
 sky130_fd_sc_hd__a21bo_1 c206 (.A1(net26),
    .A2(net684),
    .B1_N(net670),
    .X(net72));
 sky130_fd_sc_hd__a21bo_2 c207 (.A1(net60),
    .A2(net691),
    .B1_N(net693),
    .X(net73));
 sky130_fd_sc_hd__mux4_2 c208 (.A0(net73),
    .A1(net680),
    .A2(net672),
    .A3(net66),
    .S0(net810),
    .S1(net51),
    .X(net74));
 sky130_fd_sc_hd__a31o_1 c209 (.A1(net52),
    .A2(net680),
    .A3(net817),
    .B1(net74),
    .X(net75));
 sky130_fd_sc_hd__a41o_1 c210 (.A1(net74),
    .A2(net632),
    .A3(net66),
    .A4(net810),
    .B1(net832),
    .X(net76));
 sky130_fd_sc_hd__a41o_2 c211 (.A1(net70),
    .A2(net782),
    .A3(net73),
    .A4(net64),
    .B1(net855),
    .X(net77));
 sky130_fd_sc_hd__a41o_1 c212 (.A1(net68),
    .A2(net708),
    .A3(net77),
    .A4(net810),
    .B1(net664),
    .X(net78));
 sky130_fd_sc_hd__a21bo_1 c213 (.A1(net70),
    .A2(net73),
    .B1_N(net846),
    .X(net79));
 sky130_fd_sc_hd__a41o_1 c214 (.A1(net72),
    .A2(net70),
    .A3(net71),
    .A4(net832),
    .B1(net846),
    .X(net733));
 sky130_fd_sc_hd__buf_1 c215 (.A(net844),
    .X(net80));
 sky130_fd_sc_hd__a41o_2 c216 (.A1(net42),
    .A2(net808),
    .A3(net80),
    .A4(net709),
    .B1(net846),
    .X(net81));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(net77),
    .A1(net808),
    .A2(net636),
    .A3(net673),
    .S0(net79),
    .S1(net895),
    .X(net82));
 sky130_fd_sc_hd__a41o_1 c218 (.A1(net58),
    .A2(net81),
    .A3(net77),
    .A4(net808),
    .B1(net79),
    .X(net83));
 sky130_fd_sc_hd__a31o_2 c219 (.A1(net80),
    .A2(net81),
    .A3(net808),
    .B1(net844),
    .X(net762));
 sky130_fd_sc_hd__a21bo_1 c220 (.A1(net72),
    .A2(net777),
    .B1_N(net774),
    .X(net787));
 sky130_fd_sc_hd__a41o_1 c221 (.A1(net641),
    .A2(net697),
    .A3(net625),
    .A4(net721),
    .B1(net722),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 c222 (.A(net841),
    .X(net85));
 sky130_fd_sc_hd__mux4_1 c223 (.A0(net838),
    .A1(net783),
    .A2(net808),
    .A3(net710),
    .S0(net72),
    .S1(net63),
    .X(net776));
 sky130_fd_sc_hd__a21bo_1 c224 (.A1(net715),
    .A2(net797),
    .B1_N(net66),
    .X(net86));
 sky130_fd_sc_hd__a21bo_2 c225 (.A1(net710),
    .A2(net681),
    .B1_N(net685),
    .X(net87));
 sky130_fd_sc_hd__a21bo_1 c226 (.A1(net85),
    .A2(net776),
    .B1_N(net64),
    .X(net88));
 sky130_fd_sc_hd__a21bo_1 c227 (.A1(net657),
    .A2(net787),
    .B1_N(net696),
    .X(net89));
 sky130_fd_sc_hd__a21bo_1 c228 (.A1(net62),
    .A2(net698),
    .B1_N(net846),
    .X(net90));
 sky130_fd_sc_hd__a21bo_1 c229 (.A1(net38),
    .A2(net711),
    .B1_N(net811),
    .X(net91));
 sky130_fd_sc_hd__a21bo_1 c230 (.A1(net90),
    .A2(net811),
    .B1_N(net68),
    .X(net765));
 sky130_fd_sc_hd__a21bo_1 c231 (.A1(net64),
    .A2(net91),
    .B1_N(net706),
    .X(net92));
 sky130_fd_sc_hd__a41o_2 c232 (.A1(net826),
    .A2(net62),
    .A3(net833),
    .A4(net713),
    .B1(net811),
    .X(net93));
 sky130_fd_sc_hd__a41o_1 c233 (.A1(net93),
    .A2(net74),
    .A3(net646),
    .A4(net811),
    .B1(net87),
    .X(net94));
 sky130_fd_sc_hd__buf_1 c234 (.A(net841),
    .X(net95));
 sky130_fd_sc_hd__a41o_1 c235 (.A1(net811),
    .A2(net87),
    .A3(net808),
    .A4(net88),
    .B1(net810),
    .X(net96));
 sky130_fd_sc_hd__mux4_1 c236 (.A0(net670),
    .A1(net713),
    .A2(net87),
    .A3(net699),
    .S0(net54),
    .S1(clknet_1_1__leaf_net799),
    .X(net97));
 sky130_fd_sc_hd__a41o_1 c237 (.A1(net712),
    .A2(net85),
    .A3(net93),
    .A4(net811),
    .B1(clknet_1_1__leaf_net799),
    .X(net786));
 sky130_fd_sc_hd__a21bo_1 c238 (.A1(net91),
    .A2(net69),
    .B1_N(net16),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 c239 (.A(net844),
    .X(net99));
 sky130_fd_sc_hd__a21bo_1 c240 (.A1(net93),
    .A2(net70),
    .B1_N(clknet_1_1__leaf_net799),
    .X(net766));
 sky130_fd_sc_hd__a41o_1 c241 (.A1(net99),
    .A2(clknet_1_0__leaf_net766),
    .A3(net697),
    .A4(net628),
    .B1(net811),
    .X(net100));
 sky130_fd_sc_hd__mux4_2 c256 (.A0(net9),
    .A1(net11),
    .A2(net673),
    .A3(net808),
    .S0(net768),
    .S1(net693),
    .X(net779));
 sky130_fd_sc_hd__mux4_1 c257 (.A0(net746),
    .A1(clknet_1_1__leaf_net97),
    .A2(net6),
    .A3(net10),
    .S0(net13),
    .S1(net846),
    .X(net800));
 sky130_fd_sc_hd__mux4_1 c258 (.A0(clknet_1_0__leaf_net97),
    .A1(net15),
    .A2(net774),
    .A3(clknet_1_0__leaf_net800),
    .S0(net783),
    .S1(net795),
    .X(net101));
 sky130_fd_sc_hd__mux4_1 c259 (.A0(net86),
    .A1(net10),
    .A2(net794),
    .A3(net867),
    .S0(clknet_1_1__leaf_net800),
    .S1(net664),
    .X(net102));
 sky130_fd_sc_hd__mux4_1 c260 (.A0(net7),
    .A1(net14),
    .A2(clknet_1_0__leaf_net786),
    .A3(net10),
    .S0(net638),
    .S1(net903),
    .X(net742));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(net684),
    .A1(net13),
    .A2(net784),
    .A3(net779),
    .S0(net846),
    .S1(net841),
    .X(net790));
 sky130_fd_sc_hd__mux4_1 c262 (.A0(net6),
    .A1(net684),
    .A2(clknet_1_1__leaf_net800),
    .A3(net709),
    .S0(net791),
    .S1(net889),
    .X(net103));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net100),
    .A1(net779),
    .A2(net7),
    .A3(clknet_1_0__leaf_net742),
    .S0(net846),
    .S1(net841),
    .X(net104));
 sky130_fd_sc_hd__xnor2_4 c264 (.A(net853),
    .B(net820),
    .Y(net105));
 sky130_fd_sc_hd__xnor2_4 c265 (.A(net625),
    .B(net783),
    .Y(net106));
 sky130_fd_sc_hd__a21bo_1 c266 (.A1(net19),
    .A2(net635),
    .B1_N(net836),
    .X(net107));
 sky130_fd_sc_hd__xnor2_4 c267 (.A(net657),
    .B(net20),
    .Y(net108));
 sky130_fd_sc_hd__xnor2_2 c268 (.A(net635),
    .B(net106),
    .Y(net109));
 sky130_fd_sc_hd__xnor2_1 c269 (.A(net106),
    .B(net777),
    .Y(net110));
 sky130_fd_sc_hd__xnor2_4 c270 (.A(net631),
    .B(net825),
    .Y(net111));
 sky130_fd_sc_hd__a21bo_4 c271 (.A1(net824),
    .A2(net20),
    .B1_N(net17),
    .X(net112));
 sky130_fd_sc_hd__a21bo_4 c272 (.A1(net690),
    .A2(net109),
    .B1_N(net824),
    .X(net113));
 sky130_fd_sc_hd__xnor2_4 c273 (.A(net113),
    .B(net819),
    .Y(net114));
 sky130_fd_sc_hd__xnor2_4 c274 (.A(net28),
    .B(net634),
    .Y(net115));
 sky130_fd_sc_hd__a21bo_4 c275 (.A1(net105),
    .A2(net113),
    .B1_N(net849),
    .X(net116));
 sky130_fd_sc_hd__xnor2_4 c276 (.A(net819),
    .B(net635),
    .Y(net117));
 sky130_fd_sc_hd__xnor2_4 c277 (.A(net819),
    .B(net116),
    .Y(net118));
 sky130_fd_sc_hd__xnor2_4 c278 (.A(net118),
    .B(net116),
    .Y(net119));
 sky130_fd_sc_hd__a31o_2 c279 (.A1(net109),
    .A2(net113),
    .A3(net112),
    .B1(net823),
    .X(net120));
 sky130_fd_sc_hd__a31o_4 c280 (.A1(net23),
    .A2(net111),
    .A3(net668),
    .B1(net112),
    .X(net121));
 sky130_fd_sc_hd__a21bo_2 c281 (.A1(net114),
    .A2(net115),
    .B1_N(net116),
    .X(net122));
 sky130_fd_sc_hd__a41o_4 c282 (.A1(net816),
    .A2(net120),
    .A3(net122),
    .A4(net637),
    .B1(net838),
    .X(net123));
 sky130_fd_sc_hd__a21bo_4 c283 (.A1(net110),
    .A2(net122),
    .B1_N(net824),
    .X(net124));
 sky130_fd_sc_hd__mux4_2 c284 (.A0(net116),
    .A1(net122),
    .A2(net106),
    .A3(net23),
    .S0(net29),
    .S1(net838),
    .X(net125));
 sky130_fd_sc_hd__mux4_2 c285 (.A0(net122),
    .A1(net124),
    .A2(net634),
    .A3(net114),
    .S0(net111),
    .S1(net113),
    .X(net738));
 sky130_fd_sc_hd__a21bo_1 c286 (.A1(net651),
    .A2(net118),
    .B1_N(net847),
    .X(net126));
 sky130_fd_sc_hd__xnor2_2 c287 (.A(net39),
    .B(net661),
    .Y(net127));
 sky130_fd_sc_hd__xnor2_2 c288 (.A(net625),
    .B(net36),
    .Y(net128));
 sky130_fd_sc_hd__a21bo_4 c289 (.A1(net34),
    .A2(net643),
    .B1_N(net826),
    .X(net129));
 sky130_fd_sc_hd__a31o_1 c290 (.A1(net626),
    .A2(net114),
    .A3(net113),
    .B1(net655),
    .X(net130));
 sky130_fd_sc_hd__a21bo_2 c291 (.A1(net129),
    .A2(net121),
    .B1_N(net825),
    .X(net763));
 sky130_fd_sc_hd__a31o_4 c292 (.A1(net654),
    .A2(net780),
    .A3(net814),
    .B1(net852),
    .X(net131));
 sky130_fd_sc_hd__xnor2_4 c293 (.A(net131),
    .B(net814),
    .Y(net132));
 sky130_fd_sc_hd__mux4_2 c294 (.A0(net125),
    .A1(net626),
    .A2(net851),
    .A3(net847),
    .S0(net777),
    .S1(net129),
    .X(net133));
 sky130_fd_sc_hd__a31o_4 c295 (.A1(net133),
    .A2(net129),
    .A3(net638),
    .B1(net131),
    .X(net134));
 sky130_fd_sc_hd__a21bo_4 c296 (.A1(net629),
    .A2(net134),
    .B1_N(net819),
    .X(net135));
 sky130_fd_sc_hd__mux4_2 c297 (.A0(net637),
    .A1(net119),
    .A2(net33),
    .A3(net135),
    .S0(net133),
    .S1(net824),
    .X(net136));
 sky130_fd_sc_hd__mux4_2 c298 (.A0(net127),
    .A1(net23),
    .A2(net132),
    .A3(net819),
    .S0(net44),
    .S1(net829),
    .X(net137));
 sky130_fd_sc_hd__a21bo_4 c299 (.A1(net136),
    .A2(net640),
    .B1_N(net134),
    .X(net138));
 sky130_fd_sc_hd__a21bo_4 c300 (.A1(net131),
    .A2(net136),
    .B1_N(net642),
    .X(net139));
 sky130_fd_sc_hd__a21bo_1 c301 (.A1(net118),
    .A2(net129),
    .B1_N(net139),
    .X(net140));
 sky130_fd_sc_hd__a21bo_4 c302 (.A1(net139),
    .A2(net133),
    .B1_N(net138),
    .X(net141));
 sky130_fd_sc_hd__mux4_2 c303 (.A0(net138),
    .A1(net639),
    .A2(net140),
    .A3(net119),
    .S0(net690),
    .S1(net761),
    .X(net142));
 sky130_fd_sc_hd__a41o_2 c304 (.A1(net653),
    .A2(net135),
    .A3(net138),
    .A4(net814),
    .B1(net825),
    .X(net735));
 sky130_fd_sc_hd__mux4_2 c305 (.A0(net141),
    .A1(net128),
    .A2(net113),
    .A3(net122),
    .S0(net130),
    .S1(net814),
    .X(net143));
 sky130_fd_sc_hd__a21bo_4 c306 (.A1(net127),
    .A2(net121),
    .B1_N(net140),
    .X(net757));
 sky130_fd_sc_hd__a21bo_1 c307 (.A1(net143),
    .A2(net636),
    .B1_N(net757),
    .X(net144));
 sky130_fd_sc_hd__a21bo_2 c308 (.A1(net675),
    .A2(net658),
    .B1_N(net832),
    .X(net145));
 sky130_fd_sc_hd__a21bo_1 c309 (.A1(net23),
    .A2(net780),
    .B1_N(net804),
    .X(net146));
 sky130_fd_sc_hd__a21bo_4 c310 (.A1(net48),
    .A2(net33),
    .B1_N(net814),
    .X(net770));
 sky130_fd_sc_hd__a31o_2 c311 (.A1(net34),
    .A2(net126),
    .A3(net51),
    .B1(net904),
    .X(net147));
 sky130_fd_sc_hd__a21bo_1 c312 (.A1(net146),
    .A2(net48),
    .B1_N(net54),
    .X(net148));
 sky130_fd_sc_hd__a31o_1 c313 (.A1(net128),
    .A2(net896),
    .A3(net112),
    .B1(net126),
    .X(net149));
 sky130_fd_sc_hd__a21bo_2 c314 (.A1(net666),
    .A2(net665),
    .B1_N(net838),
    .X(net150));
 sky130_fd_sc_hd__a21bo_4 c315 (.A1(net848),
    .A2(net896),
    .B1_N(net56),
    .X(net151));
 sky130_fd_sc_hd__a21bo_1 c316 (.A1(net33),
    .A2(net63),
    .B1_N(net27),
    .X(net152));
 sky130_fd_sc_hd__a41o_2 c317 (.A1(net36),
    .A2(net145),
    .A3(net770),
    .A4(net839),
    .B1(net150),
    .X(net153));
 sky130_fd_sc_hd__a41o_1 c318 (.A1(net669),
    .A2(net112),
    .A3(net153),
    .A4(net138),
    .B1(net151),
    .X(net154));
 sky130_fd_sc_hd__mux4_2 c319 (.A0(net122),
    .A1(net643),
    .A2(net152),
    .A3(net145),
    .S0(net41),
    .S1(net153),
    .X(net155));
 sky130_fd_sc_hd__a21bo_1 c320 (.A1(net154),
    .A2(net48),
    .B1_N(net128),
    .X(net156));
 sky130_fd_sc_hd__a41o_1 c321 (.A1(net146),
    .A2(net155),
    .A3(net816),
    .A4(net128),
    .B1(net151),
    .X(net157));
 sky130_fd_sc_hd__mux4_2 c322 (.A0(net148),
    .A1(net51),
    .A2(net153),
    .A3(net824),
    .S0(net650),
    .S1(net831),
    .X(net158));
 sky130_fd_sc_hd__mux4_1 c323 (.A0(net138),
    .A1(net152),
    .A2(net149),
    .A3(net61),
    .S0(net833),
    .S1(clknet_1_1__leaf_net799),
    .X(net159));
 sky130_fd_sc_hd__a41o_1 c324 (.A1(net41),
    .A2(clknet_1_0__leaf_net159),
    .A3(net156),
    .A4(net674),
    .B1(net814),
    .X(net160));
 sky130_fd_sc_hd__a41o_1 c325 (.A1(net154),
    .A2(net61),
    .A3(net782),
    .A4(net770),
    .B1(clknet_1_1__leaf_net799),
    .X(net161));
 sky130_fd_sc_hd__a31o_1 c326 (.A1(net158),
    .A2(net153),
    .A3(net780),
    .B1(clknet_1_0__leaf_net799),
    .X(net162));
 sky130_fd_sc_hd__buf_2 c327 (.A(net846),
    .X(net749));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(net126),
    .A1(clknet_1_1__leaf_net161),
    .A2(net158),
    .A3(net642),
    .S0(clknet_1_1__leaf_net162),
    .S1(net770),
    .X(net163));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(clknet_1_0__leaf_net159),
    .A1(net857),
    .A2(net864),
    .A3(clknet_1_1__leaf_net162),
    .S0(clknet_1_1__leaf_net161),
    .S1(net129),
    .X(net164));
 sky130_fd_sc_hd__a41o_1 c330 (.A1(net79),
    .A2(clknet_1_1__leaf_net159),
    .A3(net804),
    .A4(net833),
    .B1(net808),
    .X(net165));
 sky130_fd_sc_hd__a21bo_1 c331 (.A1(net682),
    .A2(net821),
    .B1_N(clknet_1_1__leaf_net799),
    .X(net166));
 sky130_fd_sc_hd__a21bo_1 c332 (.A1(net80),
    .A2(net66),
    .B1_N(net821),
    .X(net167));
 sky130_fd_sc_hd__a21bo_1 c333 (.A1(clknet_1_1__leaf_net166),
    .A2(net770),
    .B1_N(net757),
    .X(net769));
 sky130_fd_sc_hd__a31o_1 c334 (.A1(net687),
    .A2(net141),
    .A3(net673),
    .B1(net821),
    .X(net168));
 sky130_fd_sc_hd__a41o_2 c335 (.A1(net780),
    .A2(net813),
    .A3(net679),
    .A4(net890),
    .B1(net846),
    .X(net169));
 sky130_fd_sc_hd__a41o_2 c336 (.A1(net658),
    .A2(net61),
    .A3(net640),
    .A4(net817),
    .B1(net49),
    .X(net755));
 sky130_fd_sc_hd__a21bo_1 c337 (.A1(net686),
    .A2(net636),
    .B1_N(net654),
    .X(net170));
 sky130_fd_sc_hd__buf_1 c338 (.A(net844),
    .X(net171));
 sky130_fd_sc_hd__a21bo_1 c339 (.A1(net635),
    .A2(net668),
    .B1_N(net71),
    .X(net773));
 sky130_fd_sc_hd__buf_1 c340 (.A(net845),
    .X(net172));
 sky130_fd_sc_hd__a31o_4 c341 (.A1(net171),
    .A2(net115),
    .A3(net167),
    .B1(net827),
    .X(net173));
 sky130_fd_sc_hd__mux4_1 c342 (.A0(net168),
    .A1(clknet_1_0__leaf_net769),
    .A2(net155),
    .A3(clknet_1_0__leaf_net166),
    .S0(net856),
    .S1(net572),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_2 c343 (.A(net572),
    .X(net754));
 sky130_fd_sc_hd__a41o_1 c344 (.A1(net172),
    .A2(net168),
    .A3(net679),
    .A4(net45),
    .B1(net687),
    .X(net175));
 sky130_fd_sc_hd__mux4_1 c345 (.A0(net890),
    .A1(net693),
    .A2(net145),
    .A3(net839),
    .S0(net827),
    .S1(net845),
    .X(net176));
 sky130_fd_sc_hd__a21bo_1 c346 (.A1(net176),
    .A2(net172),
    .B1_N(net175),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 c347 (.A0(net754),
    .A1(net172),
    .A2(net173),
    .A3(net875),
    .S0(net845),
    .S1(clknet_1_1__leaf_net799),
    .X(net178));
 sky130_fd_sc_hd__a31o_1 c348 (.A1(net175),
    .A2(net177),
    .A3(net845),
    .B1(clknet_1_1__leaf_net799),
    .X(net179));
 sky130_fd_sc_hd__a41o_1 c349 (.A1(net177),
    .A2(net773),
    .A3(net176),
    .A4(net172),
    .B1(net821),
    .X(net180));
 sky130_fd_sc_hd__a41o_1 c350 (.A1(clknet_1_1__leaf_net179),
    .A2(clknet_1_1__leaf_net178),
    .A3(net696),
    .A4(net180),
    .B1(net845),
    .X(net181));
 sky130_fd_sc_hd__a41o_4 c351 (.A1(clknet_1_0__leaf_net179),
    .A2(net760),
    .A3(net171),
    .A4(net846),
    .X(net748));
 sky130_fd_sc_hd__a21bo_1 c352 (.A1(net706),
    .A2(net690),
    .B1_N(net821),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_1 c353 (.A(net604),
    .X(net183));
 sky130_fd_sc_hd__a41o_1 c354 (.A1(net647),
    .A2(net717),
    .A3(net180),
    .A4(net706),
    .B1(net839),
    .X(net184));
 sky130_fd_sc_hd__mux4_2 c355 (.A0(net115),
    .A1(net692),
    .A2(net812),
    .A3(net778),
    .S0(net708),
    .S1(net734),
    .X(net185));
 sky130_fd_sc_hd__a41o_1 c356 (.A1(net180),
    .A2(net673),
    .A3(net857),
    .A4(net721),
    .B1(net744),
    .X(net186));
 sky130_fd_sc_hd__mux4_2 c357 (.A0(net87),
    .A1(net770),
    .A2(net762),
    .A3(net185),
    .S0(net153),
    .S1(net681),
    .X(net187));
 sky130_fd_sc_hd__a41o_1 c358 (.A1(net662),
    .A2(net185),
    .A3(net848),
    .A4(net151),
    .B1(net814),
    .X(net188));
 sky130_fd_sc_hd__a41o_1 c359 (.A1(net173),
    .A2(net810),
    .A3(net188),
    .A4(net713),
    .B1(net651),
    .X(net189));
 sky130_fd_sc_hd__a41o_1 c360 (.A1(net5),
    .A2(net690),
    .A3(net47),
    .A4(net641),
    .B1(net839),
    .X(net190));
 sky130_fd_sc_hd__a31o_1 c361 (.A1(net654),
    .A2(net702),
    .A3(net699),
    .B1(net848),
    .X(net191));
 sky130_fd_sc_hd__a31o_1 c362 (.A1(net113),
    .A2(net811),
    .A3(net185),
    .B1(net706),
    .X(net192));
 sky130_fd_sc_hd__a21bo_1 c363 (.A1(net696),
    .A2(net141),
    .B1_N(net191),
    .X(net193));
 sky130_fd_sc_hd__a31o_2 c364 (.A1(net61),
    .A2(net839),
    .A3(net190),
    .B1(net87),
    .X(net194));
 sky130_fd_sc_hd__a21bo_1 c365 (.A1(net3),
    .A2(net112),
    .B1_N(net170),
    .X(net195));
 sky130_fd_sc_hd__mux4_1 c366 (.A0(net188),
    .A1(net115),
    .A2(net783),
    .A3(net173),
    .S0(net4),
    .S1(net93),
    .X(net196));
 sky130_fd_sc_hd__mux4_2 c367 (.A0(net190),
    .A1(net147),
    .A2(net196),
    .A3(net631),
    .S0(net193),
    .S1(net713),
    .X(net197));
 sky130_fd_sc_hd__a21bo_1 c368 (.A1(net193),
    .A2(net696),
    .B1_N(clknet_1_1__leaf_net799),
    .X(net198));
 sky130_fd_sc_hd__a31o_1 c369 (.A1(net63),
    .A2(net713),
    .A3(net763),
    .B1(net638),
    .X(net750));
 sky130_fd_sc_hd__a21bo_1 c370 (.A1(net697),
    .A2(net45),
    .B1_N(clknet_1_1__leaf_net198),
    .X(net199));
 sky130_fd_sc_hd__a31o_1 c371 (.A1(net153),
    .A2(clknet_1_1__leaf_net199),
    .A3(net68),
    .B1(net844),
    .X(net200));
 sky130_fd_sc_hd__a31o_2 c372 (.A1(net170),
    .A2(net4),
    .A3(net3),
    .B1(net195),
    .X(net201));
 sky130_fd_sc_hd__a41o_1 c373 (.A1(net195),
    .A2(net817),
    .A3(clknet_1_0__leaf_net199),
    .A4(clknet_1_0__leaf_net200),
    .B1(net201),
    .X(net202));
 sky130_fd_sc_hd__xnor2_2 c396 (.A(net29),
    .B(net816),
    .Y(net203));
 sky130_fd_sc_hd__xnor2_4 c397 (.A(net628),
    .B(net120),
    .Y(net204));
 sky130_fd_sc_hd__a21bo_1 c398 (.A1(net19),
    .A2(net809),
    .B1_N(net125),
    .X(net205));
 sky130_fd_sc_hd__xnor2_2 c399 (.A(net824),
    .B(net116),
    .Y(net206));
 sky130_fd_sc_hd__a21bo_1 c400 (.A1(net204),
    .A2(net105),
    .B1_N(net120),
    .X(net207));
 sky130_fd_sc_hd__xnor2_2 c401 (.A(net820),
    .B(net631),
    .Y(net208));
 sky130_fd_sc_hd__a41o_2 c402 (.A1(net818),
    .A2(net116),
    .A3(net29),
    .A4(net626),
    .B1(net204),
    .X(net767));
 sky130_fd_sc_hd__xnor2_2 c403 (.A(net783),
    .B(net836),
    .Y(net209));
 sky130_fd_sc_hd__xnor2_2 c404 (.A(net112),
    .B(net28),
    .Y(net210));
 sky130_fd_sc_hd__a41o_4 c405 (.A1(net28),
    .A2(net208),
    .A3(net105),
    .A4(net809),
    .B1(net124),
    .X(net211));
 sky130_fd_sc_hd__a21bo_2 c406 (.A1(net207),
    .A2(net206),
    .B1_N(net809),
    .X(net212));
 sky130_fd_sc_hd__a21bo_2 c407 (.A1(net209),
    .A2(net111),
    .B1_N(net767),
    .X(net213));
 sky130_fd_sc_hd__a21bo_1 c408 (.A1(net212),
    .A2(net637),
    .B1_N(net213),
    .X(net214));
 sky130_fd_sc_hd__xnor2_4 c409 (.A(net211),
    .B(net809),
    .Y(net215));
 sky130_fd_sc_hd__mux4_2 c410 (.A0(net109),
    .A1(net628),
    .A2(net112),
    .A3(net211),
    .S0(net838),
    .S1(net809),
    .X(net216));
 sky130_fd_sc_hd__mux4_2 c411 (.A0(net631),
    .A1(net820),
    .A2(net206),
    .A3(net213),
    .S0(net824),
    .S1(net116),
    .X(net217));
 sky130_fd_sc_hd__mux4_1 c412 (.A0(net210),
    .A1(net679),
    .A2(net213),
    .A3(net809),
    .S0(net123),
    .S1(net114),
    .X(net727));
 sky130_fd_sc_hd__a21bo_1 c413 (.A1(net120),
    .A2(net809),
    .B1_N(net213),
    .X(net218));
 sky130_fd_sc_hd__a21bo_1 c414 (.A1(net217),
    .A2(net19),
    .B1_N(net211),
    .X(net219));
 sky130_fd_sc_hd__a21bo_2 c415 (.A1(net213),
    .A2(net210),
    .B1_N(net214),
    .X(net220));
 sky130_fd_sc_hd__a21bo_1 c416 (.A1(net106),
    .A2(net220),
    .B1_N(net219),
    .X(net221));
 sky130_fd_sc_hd__mux4_2 c417 (.A0(net214),
    .A1(net109),
    .A2(net809),
    .A3(net221),
    .S0(net220),
    .S1(net211),
    .X(net222));
 sky130_fd_sc_hd__a21bo_1 c418 (.A1(net134),
    .A2(net135),
    .B1_N(net825),
    .X(net223));
 sky130_fd_sc_hd__a31o_2 c419 (.A1(net908),
    .A2(net137),
    .A3(net44),
    .B1(net124),
    .X(net224));
 sky130_fd_sc_hd__mux4_2 c420 (.A0(net628),
    .A1(net123),
    .A2(net144),
    .A3(net820),
    .S0(net807),
    .S1(net39),
    .X(net225));
 sky130_fd_sc_hd__a31o_1 c421 (.A1(net636),
    .A2(net127),
    .A3(net668),
    .B1(net829),
    .X(net226));
 sky130_fd_sc_hd__a21bo_2 c422 (.A1(net226),
    .A2(net205),
    .B1_N(net829),
    .X(net227));
 sky130_fd_sc_hd__a21bo_4 c423 (.A1(net809),
    .A2(net143),
    .B1_N(net131),
    .X(net228));
 sky130_fd_sc_hd__a31o_2 c424 (.A1(net144),
    .A2(net44),
    .A3(net656),
    .B1(net223),
    .X(net229));
 sky130_fd_sc_hd__a21bo_1 c425 (.A1(net223),
    .A2(net222),
    .B1_N(net208),
    .X(net230));
 sky130_fd_sc_hd__a21bo_1 c426 (.A1(net44),
    .A2(net651),
    .B1_N(net127),
    .X(net231));
 sky130_fd_sc_hd__a21bo_2 c427 (.A1(net690),
    .A2(net230),
    .B1_N(net229),
    .X(net232));
 sky130_fd_sc_hd__a21bo_1 c428 (.A1(net656),
    .A2(net107),
    .B1_N(net215),
    .X(net233));
 sky130_fd_sc_hd__buf_1 c429 (.A(net569),
    .X(net234));
 sky130_fd_sc_hd__a31o_1 c430 (.A1(net232),
    .A2(net135),
    .A3(net123),
    .B1(net233),
    .X(net235));
 sky130_fd_sc_hd__a21bo_2 c431 (.A1(net234),
    .A2(net230),
    .B1_N(net130),
    .X(net236));
 sky130_fd_sc_hd__a21bo_1 c432 (.A1(net659),
    .A2(net125),
    .B1_N(net227),
    .X(net237));
 sky130_fd_sc_hd__a21bo_1 c433 (.A1(net32),
    .A2(net881),
    .B1_N(net211),
    .X(net238));
 sky130_fd_sc_hd__a21bo_2 c434 (.A1(net20),
    .A2(net134),
    .B1_N(net626),
    .X(net239));
 sky130_fd_sc_hd__mux4_1 c435 (.A0(net227),
    .A1(net212),
    .A2(net220),
    .A3(net229),
    .S0(net234),
    .S1(net237),
    .X(net240));
 sky130_fd_sc_hd__a31o_1 c436 (.A1(net130),
    .A2(net637),
    .A3(net240),
    .B1(net238),
    .X(net241));
 sky130_fd_sc_hd__a31o_1 c437 (.A1(net231),
    .A2(net205),
    .A3(net203),
    .B1(net42),
    .X(net242));
 sky130_fd_sc_hd__a21bo_1 c438 (.A1(net144),
    .A2(net731),
    .B1_N(net843),
    .X(net243));
 sky130_fd_sc_hd__a31o_1 c439 (.A1(net140),
    .A2(net243),
    .A3(net809),
    .B1(net842),
    .X(net244));
 sky130_fd_sc_hd__a41o_1 c440 (.A1(net231),
    .A2(net656),
    .A3(net829),
    .A4(net119),
    .B1(net242),
    .X(net245));
 sky130_fd_sc_hd__a21bo_1 c441 (.A1(net641),
    .A2(net42),
    .B1_N(net814),
    .X(net246));
 sky130_fd_sc_hd__a21bo_1 c442 (.A1(net154),
    .A2(net150),
    .B1_N(net59),
    .X(net247));
 sky130_fd_sc_hd__dlymetal6s2s_1 c443 (.A(net843),
    .X(net248));
 sky130_fd_sc_hd__a41o_2 c444 (.A1(net226),
    .A2(net671),
    .A3(net248),
    .A4(net142),
    .B1(net42),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_1 c445 (.A(net843),
    .X(net250));
 sky130_fd_sc_hd__a21bo_2 c446 (.A1(net222),
    .A2(net123),
    .B1_N(net767),
    .X(net737));
 sky130_fd_sc_hd__a21bo_1 c447 (.A1(net685),
    .A2(net672),
    .B1_N(net683),
    .X(net251));
 sky130_fd_sc_hd__a21bo_1 c448 (.A1(net45),
    .A2(net236),
    .B1_N(net897),
    .X(net252));
 sky130_fd_sc_hd__mux4_1 c449 (.A0(net240),
    .A1(net239),
    .A2(net150),
    .A3(net59),
    .S0(net151),
    .S1(clknet_1_0__leaf_net799),
    .X(net253));
 sky130_fd_sc_hd__a21bo_1 c450 (.A1(net246),
    .A2(net149),
    .B1_N(net220),
    .X(net254));
 sky130_fd_sc_hd__a41o_1 c451 (.A1(net248),
    .A2(net247),
    .A3(net683),
    .A4(net252),
    .B1(clknet_1_0__leaf_net799),
    .X(net255));
 sky130_fd_sc_hd__a41o_1 c452 (.A1(net659),
    .A2(net248),
    .A3(net814),
    .A4(net896),
    .B1(clknet_1_1__leaf_net162),
    .X(net256));
 sky130_fd_sc_hd__a21bo_1 c453 (.A1(net249),
    .A2(net142),
    .B1_N(net132),
    .X(net257));
 sky130_fd_sc_hd__mux4_1 c454 (.A0(net251),
    .A1(net247),
    .A2(net257),
    .A3(net245),
    .S0(net151),
    .S1(net603),
    .X(net258));
 sky130_fd_sc_hd__mux4_2 c455 (.A0(net245),
    .A1(net56),
    .A2(net151),
    .A3(net668),
    .S0(net878),
    .S1(net842),
    .X(net259));
 sky130_fd_sc_hd__a31o_2 c456 (.A1(net257),
    .A2(net251),
    .A3(net259),
    .B1(net57),
    .X(net260));
 sky130_fd_sc_hd__mux4_2 c457 (.A0(net147),
    .A1(net40),
    .A2(net47),
    .A3(net757),
    .S0(net259),
    .S1(net603),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_2 c458 (.A(net604),
    .X(net262));
 sky130_fd_sc_hd__a21bo_1 c459 (.A1(net262),
    .A2(net664),
    .B1_N(net237),
    .X(net263));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net259),
    .A1(net260),
    .A2(net246),
    .A3(net263),
    .S0(net261),
    .S1(net770),
    .X(net264));
 sky130_fd_sc_hd__mux4_2 c461 (.A0(net263),
    .A1(net805),
    .A2(net156),
    .A3(net261),
    .S0(net249),
    .S1(net248),
    .X(net265));
 sky130_fd_sc_hd__a31o_1 c462 (.A1(net239),
    .A2(net245),
    .A3(net254),
    .B1(net834),
    .X(net266));
 sky130_fd_sc_hd__a41o_1 c463 (.A1(net142),
    .A2(net262),
    .A3(net770),
    .A4(net681),
    .B1(net603),
    .X(net267));
 sky130_fd_sc_hd__a41o_1 c464 (.A1(net650),
    .A2(net705),
    .A3(net67),
    .A4(net734),
    .B1(clknet_1_0__leaf_net799),
    .X(net268));
 sky130_fd_sc_hd__a41o_1 c465 (.A1(net51),
    .A2(net220),
    .A3(clknet_1_1__leaf_net162),
    .A4(clknet_1_1__leaf_net268),
    .B1(net232),
    .X(net269));
 sky130_fd_sc_hd__a41o_2 c466 (.A1(net167),
    .A2(net262),
    .A3(net875),
    .A4(net145),
    .B1(net734),
    .X(net270));
 sky130_fd_sc_hd__a41o_2 c467 (.A1(net267),
    .A2(net805),
    .A3(net65),
    .A4(net707),
    .B1(net603),
    .X(net271));
 sky130_fd_sc_hd__mux4_1 c468 (.A0(net67),
    .A1(net250),
    .A2(net770),
    .A3(net810),
    .S0(net847),
    .S1(net830),
    .X(net272));
 sky130_fd_sc_hd__mux4_1 c469 (.A0(net149),
    .A1(net815),
    .A2(net683),
    .A3(net229),
    .S0(net239),
    .S1(net270),
    .X(net273));
 sky130_fd_sc_hd__a31o_1 c470 (.A1(net150),
    .A2(net271),
    .A3(net262),
    .B1(net68),
    .X(net274));
 sky130_fd_sc_hd__mux4_1 c471 (.A0(net208),
    .A1(net762),
    .A2(net749),
    .A3(net150),
    .S0(net851),
    .S1(net830),
    .X(net275));
 sky130_fd_sc_hd__a41o_1 c472 (.A1(net229),
    .A2(net271),
    .A3(net254),
    .A4(net677),
    .B1(clknet_1_1__leaf_net178),
    .X(net276));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(net156),
    .A1(net51),
    .A2(net67),
    .A3(clknet_1_0__leaf_net178),
    .S0(net805),
    .S1(net169),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 c474 (.A0(net254),
    .A1(net628),
    .A2(net54),
    .A3(net810),
    .S0(net151),
    .S1(net679),
    .X(net278));
 sky130_fd_sc_hd__mux4_1 c475 (.A0(net119),
    .A1(net808),
    .A2(net757),
    .A3(net272),
    .S0(net229),
    .S1(net843),
    .X(net279));
 sky130_fd_sc_hd__a41o_1 c476 (.A1(net279),
    .A2(net49),
    .A3(net273),
    .A4(net757),
    .B1(net265),
    .X(net280));
 sky130_fd_sc_hd__a41o_1 c477 (.A1(net707),
    .A2(net229),
    .A3(net642),
    .A4(net844),
    .B1(net843),
    .X(net736));
 sky130_fd_sc_hd__a41o_1 c478 (.A1(net688),
    .A2(net677),
    .A3(net707),
    .A4(clknet_1_1__leaf_net277),
    .B1(net834),
    .X(net281));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(clknet_1_1__leaf_net281),
    .A1(net112),
    .A2(net42),
    .A3(net239),
    .S0(net66),
    .S1(net271),
    .X(net282));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net705),
    .A1(net274),
    .A2(net271),
    .A3(net81),
    .S0(clknet_1_0__leaf_net281),
    .S1(net753),
    .X(net283));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(clknet_1_0__leaf_net277),
    .A1(net278),
    .A2(net252),
    .A3(net274),
    .S0(net271),
    .S1(clknet_1_0__leaf_net281),
    .X(net284));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(net691),
    .A1(net736),
    .A2(clknet_1_0__leaf_net282),
    .A3(net709),
    .S0(net592),
    .S1(net603),
    .X(net285));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net250),
    .A1(net37),
    .A2(net767),
    .A3(net77),
    .S0(net279),
    .S1(net822),
    .X(net286));
 sky130_fd_sc_hd__a41o_1 c484 (.A1(net270),
    .A2(clknet_1_1__leaf_net200),
    .A3(net47),
    .A4(net685),
    .B1(net804),
    .X(net287));
 sky130_fd_sc_hd__mux4_1 c485 (.A0(net4),
    .A1(net713),
    .A2(net755),
    .A3(net722),
    .S0(net738),
    .S1(net629),
    .X(net288));
 sky130_fd_sc_hd__mux4_2 c486 (.A0(net700),
    .A1(net642),
    .A2(net817),
    .A3(net639),
    .S0(net804),
    .S1(net603),
    .X(net764));
 sky130_fd_sc_hd__mux4_2 c487 (.A0(net220),
    .A1(net57),
    .A2(net699),
    .A3(net814),
    .S0(net818),
    .S1(clknet_1_0__leaf_net799),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 c488 (.A0(net95),
    .A1(net90),
    .A2(net189),
    .A3(net220),
    .S0(net693),
    .S1(net812),
    .X(net290));
 sky130_fd_sc_hd__mux4_1 c489 (.A0(net151),
    .A1(net260),
    .A2(net201),
    .A3(net749),
    .S0(net817),
    .S1(net649),
    .X(net291));
 sky130_fd_sc_hd__mux4_1 c490 (.A0(net721),
    .A1(net631),
    .A2(net247),
    .A3(clknet_1_1__leaf_net289),
    .S0(net811),
    .S1(net821),
    .X(net292));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(net147),
    .A1(net66),
    .A2(net758),
    .A3(net65),
    .S0(net677),
    .S1(clknet_1_0__leaf_net766),
    .X(net293));
 sky130_fd_sc_hd__mux4_1 c492 (.A0(net47),
    .A1(net65),
    .A2(net674),
    .A3(net754),
    .S0(net762),
    .S1(net66),
    .X(net745));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(clknet_1_1__leaf_net282),
    .A1(net764),
    .A2(net765),
    .A3(net690),
    .S0(net757),
    .S1(net746),
    .X(net294));
 sky130_fd_sc_hd__mux4_2 c494 (.A0(clknet_1_0__leaf_net289),
    .A1(net183),
    .A2(net270),
    .A3(net114),
    .S0(net151),
    .S1(clknet_1_0__leaf_net799),
    .X(net295));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(net896),
    .A1(net49),
    .A2(net270),
    .A3(net827),
    .S0(net592),
    .S1(net612),
    .X(net296));
 sky130_fd_sc_hd__a41o_1 c496 (.A1(net649),
    .A2(net746),
    .A3(clknet_1_1__leaf_net276),
    .A4(clknet_1_0__leaf_net769),
    .B1(net613),
    .X(net297));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net639),
    .A1(net886),
    .A2(net224),
    .A3(net201),
    .S0(net783),
    .S1(net804),
    .X(net298));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(net290),
    .A1(net653),
    .A2(net192),
    .A3(net270),
    .S0(net734),
    .S1(net821),
    .X(net299));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(net677),
    .A1(net298),
    .A2(net270),
    .A3(net750),
    .S0(clknet_1_1__leaf_net295),
    .S1(net834),
    .X(net300));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(net292),
    .A1(net764),
    .A2(net98),
    .A3(net744),
    .S0(net201),
    .S1(net841),
    .X(net301));
 sky130_fd_sc_hd__mux4_2 c501 (.A0(net119),
    .A1(net296),
    .A2(net755),
    .A3(net811),
    .S0(net851),
    .S1(net865),
    .X(net302));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(net56),
    .A1(net754),
    .A2(clknet_1_1__leaf_net300),
    .A3(clknet_1_1__leaf_net198),
    .S0(net173),
    .S1(net600),
    .X(net303));
 sky130_fd_sc_hd__a41o_1 c503 (.A1(net183),
    .A2(clknet_1_0__leaf_net300),
    .A3(clknet_1_0__leaf_net301),
    .A4(net194),
    .B1(net821),
    .X(net304));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net674),
    .A1(net626),
    .A2(clknet_1_1__leaf_net301),
    .A3(net672),
    .S0(net649),
    .S1(clknet_1_1__leaf_net289),
    .X(net305));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(net299),
    .A1(net717),
    .A2(clknet_1_1__leaf_net305),
    .A3(net725),
    .S0(clknet_1_1__leaf_net198),
    .S1(net600),
    .X(net306));
 sky130_fd_sc_hd__a21bo_4 c528 (.A1(net634),
    .A2(net111),
    .B1_N(net211),
    .X(net307));
 sky130_fd_sc_hd__xnor2_2 c529 (.A(net121),
    .B(net111),
    .Y(net308));
 sky130_fd_sc_hd__xnor2_4 c530 (.A(net852),
    .B(net307),
    .Y(net309));
 sky130_fd_sc_hd__xnor2_4 c531 (.A(net836),
    .B(net637),
    .Y(net310));
 sky130_fd_sc_hd__a31o_4 c532 (.A1(net211),
    .A2(net852),
    .A3(net210),
    .B1(net310),
    .X(net311));
 sky130_fd_sc_hd__mux4_2 c533 (.A0(net213),
    .A1(net309),
    .A2(net307),
    .A3(net121),
    .S0(net634),
    .S1(net806),
    .X(net312));
 sky130_fd_sc_hd__xnor2_2 c534 (.A(net309),
    .B(net218),
    .Y(net313));
 sky130_fd_sc_hd__xnor2_4 c535 (.A(net312),
    .B(net310),
    .Y(net314));
 sky130_fd_sc_hd__xnor2_4 c536 (.A(net204),
    .B(net312),
    .Y(net315));
 sky130_fd_sc_hd__a31o_4 c537 (.A1(net761),
    .A2(net221),
    .A3(net21),
    .B1(net828),
    .X(net316));
 sky130_fd_sc_hd__a31o_4 c538 (.A1(net206),
    .A2(net21),
    .A3(net313),
    .B1(net312),
    .X(net317));
 sky130_fd_sc_hd__xnor2_4 c539 (.A(net838),
    .B(net309),
    .Y(net318));
 sky130_fd_sc_hd__xnor2_4 c540 (.A(net316),
    .B(net315),
    .Y(net726));
 sky130_fd_sc_hd__a21bo_1 c541 (.A1(net316),
    .A2(net207),
    .B1_N(net206),
    .X(net319));
 sky130_fd_sc_hd__xnor2_1 c542 (.A(net105),
    .B(net124),
    .Y(net320));
 sky130_fd_sc_hd__a21bo_1 c543 (.A1(net317),
    .A2(net314),
    .B1_N(net806),
    .X(net321));
 sky130_fd_sc_hd__mux4_2 c544 (.A0(net319),
    .A1(net307),
    .A2(net318),
    .A3(net816),
    .S0(net311),
    .S1(net668),
    .X(net322));
 sky130_fd_sc_hd__a31o_1 c545 (.A1(net314),
    .A2(net312),
    .A3(net123),
    .B1(net29),
    .X(net323));
 sky130_fd_sc_hd__a31o_1 c546 (.A1(net207),
    .A2(net679),
    .A3(net320),
    .B1(net313),
    .X(net324));
 sky130_fd_sc_hd__mux4_2 c547 (.A0(net321),
    .A1(net313),
    .A2(net324),
    .A3(net209),
    .S0(net316),
    .S1(net806),
    .X(net325));
 sky130_fd_sc_hd__a41o_2 c548 (.A1(net111),
    .A2(net323),
    .A3(net325),
    .A4(net215),
    .B1(net314),
    .X(net326));
 sky130_fd_sc_hd__a31o_1 c549 (.A1(net326),
    .A2(net316),
    .A3(net213),
    .B1(net325),
    .X(net327));
 sky130_fd_sc_hd__a41o_4 c550 (.A1(net133),
    .A2(net315),
    .A3(net314),
    .A4(net625),
    .B1(net602),
    .X(net723));
 sky130_fd_sc_hd__a41o_2 c551 (.A1(net39),
    .A2(net325),
    .A3(net138),
    .A4(net322),
    .B1(net723),
    .X(net752));
 sky130_fd_sc_hd__a31o_1 c552 (.A1(net661),
    .A2(net30),
    .A3(net317),
    .B1(net211),
    .X(net328));
 sky130_fd_sc_hd__a21bo_1 c553 (.A1(net328),
    .A2(net816),
    .B1_N(net890),
    .X(net329));
 sky130_fd_sc_hd__a21bo_1 c554 (.A1(net238),
    .A2(net43),
    .B1_N(net819),
    .X(net330));
 sky130_fd_sc_hd__a31o_1 c555 (.A1(net321),
    .A2(net723),
    .A3(net327),
    .B1(net138),
    .X(net331));
 sky130_fd_sc_hd__a41o_1 c556 (.A1(net135),
    .A2(net232),
    .A3(net121),
    .A4(net39),
    .B1(net227),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_1 c557 (.A(net562),
    .X(net333));
 sky130_fd_sc_hd__a31o_2 c558 (.A1(net333),
    .A2(net137),
    .A3(net225),
    .B1(net825),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_1 c559 (.A(net562),
    .X(net335));
 sky130_fd_sc_hd__a31o_1 c560 (.A1(net230),
    .A2(net752),
    .A3(net807),
    .B1(net825),
    .X(net336));
 sky130_fd_sc_hd__a31o_1 c561 (.A1(net335),
    .A2(net25),
    .A3(net806),
    .B1(net573),
    .X(net337));
 sky130_fd_sc_hd__a31o_1 c562 (.A1(net221),
    .A2(net336),
    .A3(net328),
    .B1(net753),
    .X(net338));
 sky130_fd_sc_hd__buf_1 c563 (.A(net569),
    .X(net339));
 sky130_fd_sc_hd__a31o_1 c564 (.A1(net339),
    .A2(net318),
    .A3(net43),
    .B1(net824),
    .X(net340));
 sky130_fd_sc_hd__mux4_2 c565 (.A0(net337),
    .A1(net314),
    .A2(net131),
    .A3(net340),
    .S0(net339),
    .S1(net660),
    .X(net341));
 sky130_fd_sc_hd__mux4_2 c566 (.A0(net203),
    .A1(net39),
    .A2(net881),
    .A3(net25),
    .S0(net819),
    .S1(net333),
    .X(net747));
 sky130_fd_sc_hd__sdfbbn_1 c567 (.CLK_N(clknet_2_0__leaf_clk),
    .D(net313),
    .RESET_B(net338),
    .SCD(net747),
    .SCE(net341),
    .SET_B(net657),
    .Q(net343),
    .Q_N(net342));
 sky130_fd_sc_hd__a31o_1 c568 (.A1(net338),
    .A2(net336),
    .A3(net804),
    .B1(net322),
    .X(net344));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(net655),
    .A1(net747),
    .A2(net330),
    .A3(net752),
    .S0(net236),
    .S1(net574),
    .X(net345));
 sky130_fd_sc_hd__a41o_2 c570 (.A1(net804),
    .A2(net329),
    .A3(net337),
    .A4(net342),
    .B1(net574),
    .X(net346));
 sky130_fd_sc_hd__mux4_1 c571 (.A0(net205),
    .A1(net338),
    .A2(net342),
    .A3(net330),
    .S0(net747),
    .S1(net574),
    .X(net347));
 sky130_fd_sc_hd__a21bo_1 c572 (.A1(net340),
    .A2(net858),
    .B1_N(net645),
    .X(net348));
 sky130_fd_sc_hd__a41o_1 c573 (.A1(net260),
    .A2(net848),
    .A3(net329),
    .A4(net222),
    .B1(net830),
    .X(net349));
 sky130_fd_sc_hd__a41o_1 c574 (.A1(net904),
    .A2(net858),
    .A3(clknet_1_0__leaf_net162),
    .A4(net807),
    .B1(net16),
    .X(net350));
 sky130_fd_sc_hd__a21bo_1 c575 (.A1(net322),
    .A2(net672),
    .B1_N(net671),
    .X(net351));
 sky130_fd_sc_hd__mux4_1 c576 (.A0(net236),
    .A1(net146),
    .A2(net737),
    .A3(net42),
    .S0(net265),
    .S1(clknet_1_0__leaf_net161),
    .X(net352));
 sky130_fd_sc_hd__a21bo_2 c577 (.A1(net251),
    .A2(net569),
    .B1_N(net743),
    .X(net353));
 sky130_fd_sc_hd__a21bo_2 c578 (.A1(net336),
    .A2(net850),
    .B1_N(net216),
    .X(net354));
 sky130_fd_sc_hd__mux4_1 c579 (.A0(net330),
    .A1(net341),
    .A2(net850),
    .A3(net679),
    .S0(net870),
    .S1(net569),
    .X(net355));
 sky130_fd_sc_hd__a21bo_1 c580 (.A1(net261),
    .A2(net657),
    .B1_N(net236),
    .X(net356));
 sky130_fd_sc_hd__a41o_1 c581 (.A1(net335),
    .A2(net904),
    .A3(net839),
    .A4(net242),
    .B1(net353),
    .X(net357));
 sky130_fd_sc_hd__a31o_1 c582 (.A1(net237),
    .A2(net357),
    .A3(net807),
    .B1(net892),
    .X(net358));
 sky130_fd_sc_hd__a21bo_1 c583 (.A1(net879),
    .A2(net341),
    .B1_N(net743),
    .X(net359));
 sky130_fd_sc_hd__mux4_1 c584 (.A0(net679),
    .A1(net660),
    .A2(net829),
    .A3(net341),
    .S0(net816),
    .S1(net353),
    .X(net360));
 sky130_fd_sc_hd__a31o_1 c585 (.A1(net132),
    .A2(net637),
    .A3(net338),
    .B1(net327),
    .X(net361));
 sky130_fd_sc_hd__a41o_1 c586 (.A1(net356),
    .A2(net358),
    .A3(net334),
    .A4(net131),
    .B1(net357),
    .X(net362));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(net360),
    .A1(net338),
    .A2(net343),
    .A3(net356),
    .S0(net650),
    .S1(net850),
    .X(net363));
 sky130_fd_sc_hd__a41o_1 c588 (.A1(net327),
    .A2(net353),
    .A3(net237),
    .A4(net336),
    .B1(clknet_1_0__leaf_net162),
    .X(net364));
 sky130_fd_sc_hd__mux4_1 c589 (.A0(clknet_1_0__leaf_net161),
    .A1(net353),
    .A2(net341),
    .A3(net354),
    .S0(net807),
    .S1(net618),
    .X(net365));
 sky130_fd_sc_hd__a21bo_1 c590 (.A1(net359),
    .A2(net318),
    .B1_N(clknet_1_0__leaf_net614),
    .X(net366));
 sky130_fd_sc_hd__a21bo_1 c591 (.A1(net366),
    .A2(net257),
    .B1_N(net359),
    .X(net367));
 sky130_fd_sc_hd__mux4_1 c592 (.A0(net324),
    .A1(net353),
    .A2(net227),
    .A3(net236),
    .S0(net597),
    .S1(net841),
    .X(net368));
 sky130_fd_sc_hd__a41o_1 c593 (.A1(net152),
    .A2(net353),
    .A3(clknet_1_1__leaf_net367),
    .A4(net312),
    .B1(net841),
    .X(net369));
 sky130_fd_sc_hd__mux4_1 c594 (.A0(net81),
    .A1(net692),
    .A2(net138),
    .A3(net341),
    .S0(net657),
    .S1(clknet_1_0__leaf_net799),
    .X(net370));
 sky130_fd_sc_hd__mux4_2 c595 (.A0(net650),
    .A1(net138),
    .A2(net737),
    .A3(net182),
    .S0(net835),
    .S1(net886),
    .X(net751));
 sky130_fd_sc_hd__mux4_1 c596 (.A0(net169),
    .A1(net129),
    .A2(net851),
    .A3(net848),
    .S0(net734),
    .S1(net604),
    .X(net371));
 sky130_fd_sc_hd__a41o_1 c597 (.A1(net645),
    .A2(net42),
    .A3(net224),
    .A4(net878),
    .B1(net822),
    .X(net372));
 sky130_fd_sc_hd__a41o_1 c598 (.A1(net271),
    .A2(net267),
    .A3(net819),
    .A4(net312),
    .B1(net839),
    .X(net373));
 sky130_fd_sc_hd__a41o_1 c599 (.A1(clknet_1_0__leaf_net268),
    .A2(net319),
    .A3(net749),
    .A4(net271),
    .B1(net667),
    .X(net374));
 sky130_fd_sc_hd__mux4_1 c600 (.A0(clknet_1_0__leaf_net178),
    .A1(net169),
    .A2(net59),
    .A3(net341),
    .S0(net597),
    .S1(net616),
    .X(net375));
 sky130_fd_sc_hd__a41o_1 c601 (.A1(clknet_1_1__leaf_net375),
    .A2(net77),
    .A3(net373),
    .A4(net351),
    .B1(net602),
    .X(net376));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(net30),
    .A1(net232),
    .A2(net307),
    .A3(net874),
    .S0(net808),
    .S1(net743),
    .X(net377));
 sky130_fd_sc_hd__a41o_1 c603 (.A1(net371),
    .A2(net326),
    .A3(net835),
    .A4(net329),
    .B1(net858),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(net679),
    .A1(net232),
    .A2(net307),
    .A3(net312),
    .S0(net372),
    .S1(net827),
    .X(net379));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net374),
    .A1(net334),
    .A2(net698),
    .A3(net351),
    .S0(net326),
    .S1(clknet_1_0__leaf_net799),
    .X(net380));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net252),
    .A1(net665),
    .A2(net815),
    .A3(net709),
    .S0(net681),
    .S1(net844),
    .X(net381));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(net685),
    .A1(net353),
    .A2(net650),
    .A3(net871),
    .S0(net573),
    .S1(net759),
    .X(net382));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net341),
    .A1(net275),
    .A2(net751),
    .A3(net850),
    .S0(net752),
    .S1(net679),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 c609 (.A0(net629),
    .A1(net382),
    .A2(net372),
    .A3(net312),
    .S0(net876),
    .S1(net743),
    .X(net384));
 sky130_fd_sc_hd__mux4_1 c610 (.A0(net325),
    .A1(net645),
    .A2(net275),
    .A3(net114),
    .S0(clknet_1_0__leaf_net255),
    .S1(net382),
    .X(net385));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net384),
    .A1(net311),
    .A2(net317),
    .A3(clknet_1_0__leaf_net375),
    .S0(clknet_1_0__leaf_net162),
    .S1(net842),
    .X(net386));
 sky130_fd_sc_hd__a41o_2 c612 (.A1(net329),
    .A2(net683),
    .A3(net738),
    .A4(net692),
    .B1(net608),
    .X(net387));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(net81),
    .A1(net709),
    .A2(net54),
    .A3(net691),
    .S0(net387),
    .S1(net608),
    .X(net388));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(net385),
    .A1(net372),
    .A2(net224),
    .A3(net387),
    .S0(net625),
    .S1(net629),
    .X(net389));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net388),
    .A1(net387),
    .A2(net114),
    .A3(net726),
    .S0(net759),
    .S1(clknet_1_1__leaf_net614),
    .X(net793));
 sky130_fd_sc_hd__mux4_2 c616 (.A0(net387),
    .A1(net189),
    .A2(net732),
    .A3(net847),
    .S0(net749),
    .S1(net821),
    .X(net739));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(net272),
    .A1(net804),
    .A2(net805),
    .A3(net629),
    .S0(net835),
    .S1(net841),
    .X(net390));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(net247),
    .A1(clknet_1_0__leaf_net305),
    .A2(net685),
    .A3(net173),
    .S0(net801),
    .S1(clknet_1_1__leaf_net799),
    .X(net391));
 sky130_fd_sc_hd__mux4_1 c619 (.A0(clknet_1_1__leaf_net295),
    .A1(net191),
    .A2(net73),
    .A3(clknet_1_1__leaf_net301),
    .S0(net834),
    .S1(net592),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net351),
    .A1(net668),
    .A2(net699),
    .A3(clknet_1_0__leaf_net198),
    .S0(net722),
    .S1(net612),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(net381),
    .A1(net348),
    .A2(net265),
    .A3(clknet_1_0__leaf_net289),
    .S0(net805),
    .S1(net844),
    .X(net394));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(net672),
    .A1(net201),
    .A2(net702),
    .A3(net847),
    .S0(net759),
    .S1(net612),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(net224),
    .A1(net394),
    .A2(net182),
    .A3(net657),
    .S0(net737),
    .S1(clknet_1_0__leaf_net793),
    .X(net396));
 sky130_fd_sc_hd__mux4_1 c624 (.A0(net196),
    .A1(net182),
    .A2(net260),
    .A3(net224),
    .S0(net608),
    .S1(net613),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net378),
    .A1(net643),
    .A2(clknet_1_0__leaf_net295),
    .A3(net667),
    .S0(net725),
    .S1(net593),
    .X(net398));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(clknet_1_0__leaf_net276),
    .A1(net395),
    .A2(net651),
    .A3(net804),
    .S0(net191),
    .S1(net822),
    .X(net399));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(net145),
    .A1(net54),
    .A2(clknet_1_1__leaf_net255),
    .A3(net625),
    .S0(net387),
    .S1(net620),
    .X(net741));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net685),
    .A1(net173),
    .A2(clknet_1_0__leaf_net295),
    .A3(net815),
    .S0(net851),
    .S1(net593),
    .X(net400));
 sky130_fd_sc_hd__a41o_1 c629 (.A1(net201),
    .A2(net851),
    .A3(net354),
    .A4(net603),
    .B1(net621),
    .X(net401));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net390),
    .A1(net197),
    .A2(net804),
    .A3(net672),
    .S0(net812),
    .S1(net816),
    .X(net402));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net114),
    .A1(clknet_1_1__leaf_net289),
    .A2(net626),
    .A3(net593),
    .S0(net801),
    .S1(net620),
    .X(net403));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net651),
    .A1(net403),
    .A2(net197),
    .A3(net54),
    .S0(net387),
    .S1(clknet_1_1__leaf_net400),
    .X(net404));
 sky130_fd_sc_hd__mux4_2 c633 (.A0(net273),
    .A1(net395),
    .A2(net723),
    .A3(net351),
    .S0(net734),
    .S1(net612),
    .X(net405));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(clknet_1_0__leaf_net198),
    .A1(net192),
    .A2(clknet_1_0__leaf_net289),
    .A3(net387),
    .S0(net801),
    .S1(net621),
    .X(net406));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net84),
    .A1(net683),
    .A2(net746),
    .A3(net759),
    .S0(net611),
    .S1(clknet_1_1__leaf_net615),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net98),
    .A1(clknet_1_0__leaf_net301),
    .A2(net668),
    .A3(net685),
    .S0(net849),
    .S1(net611),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net383),
    .A1(net408),
    .A2(net723),
    .A3(net593),
    .S0(clknet_1_1__leaf_net615),
    .S1(net621),
    .X(net409));
 sky130_fd_sc_hd__a31o_2 c660 (.A1(net309),
    .A2(net311),
    .A3(net828),
    .B1(net860),
    .X(net410));
 sky130_fd_sc_hd__a21bo_1 c661 (.A1(net218),
    .A2(net308),
    .B1_N(net322),
    .X(net411));
 sky130_fd_sc_hd__a41o_2 c662 (.A1(net217),
    .A2(net316),
    .A3(net411),
    .A4(net818),
    .B1(net807),
    .X(net412));
 sky130_fd_sc_hd__xnor2_2 c663 (.A(net214),
    .B(net323),
    .Y(net413));
 sky130_fd_sc_hd__xnor2_1 c664 (.A(net209),
    .B(net726),
    .Y(net414));
 sky130_fd_sc_hd__a21bo_2 c665 (.A1(net411),
    .A2(net219),
    .B1_N(net818),
    .X(net415));
 sky130_fd_sc_hd__a31o_1 c666 (.A1(net219),
    .A2(net887),
    .A3(net212),
    .B1(net322),
    .X(net416));
 sky130_fd_sc_hd__a21bo_1 c667 (.A1(net123),
    .A2(net308),
    .B1_N(net413),
    .X(net417));
 sky130_fd_sc_hd__a41o_1 c668 (.A1(net417),
    .A2(net410),
    .A3(net307),
    .A4(net317),
    .B1(net124),
    .X(net418));
 sky130_fd_sc_hd__a41o_1 c669 (.A1(net323),
    .A2(net413),
    .A3(net317),
    .A4(net807),
    .B1(net411),
    .X(net419));
 sky130_fd_sc_hd__a21bo_1 c670 (.A1(net210),
    .A2(net413),
    .B1_N(net847),
    .X(net420));
 sky130_fd_sc_hd__a21bo_1 c671 (.A1(net418),
    .A2(net824),
    .B1_N(net869),
    .X(net421));
 sky130_fd_sc_hd__a31o_1 c672 (.A1(net888),
    .A2(net738),
    .A3(net420),
    .B1(net862),
    .X(net422));
 sky130_fd_sc_hd__a21bo_1 c673 (.A1(net420),
    .A2(net418),
    .B1_N(net317),
    .X(net423));
 sky130_fd_sc_hd__a21bo_2 c674 (.A1(net861),
    .A2(net124),
    .B1_N(net416),
    .X(net724));
 sky130_fd_sc_hd__a21bo_2 c675 (.A1(net413),
    .A2(net724),
    .B1_N(net420),
    .X(net424));
 sky130_fd_sc_hd__a41o_1 c676 (.A1(net419),
    .A2(net861),
    .A3(net424),
    .A4(net423),
    .B1(net116),
    .X(net425));
 sky130_fd_sc_hd__sdfbbn_1 c677 (.CLK_N(clknet_2_0__leaf_clk),
    .D(net414),
    .RESET_B(net411),
    .SCD(net124),
    .SCE(net424),
    .SET_B(net418),
    .Q(net427),
    .Q_N(net426));
 sky130_fd_sc_hd__sdfbbp_1 c678 (.CLK(clknet_2_0__leaf_clk),
    .D(net116),
    .RESET_B(net308),
    .SCD(net424),
    .SCE(net415),
    .SET_B(net823),
    .Q(net429),
    .Q_N(net428));
 sky130_fd_sc_hd__a41o_1 c679 (.A1(net421),
    .A2(net894),
    .A3(net218),
    .A4(net424),
    .B1(net217),
    .X(net430));
 sky130_fd_sc_hd__a41o_1 c680 (.A1(net422),
    .A2(net424),
    .A3(net427),
    .A4(net116),
    .B1(net322),
    .X(net431));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(net424),
    .A1(net428),
    .A2(net863),
    .A3(net316),
    .S0(net543),
    .S1(net571),
    .X(net432));
 sky130_fd_sc_hd__mux4_1 c682 (.A0(net625),
    .A1(net243),
    .A2(net310),
    .A3(net657),
    .S0(net412),
    .S1(net843),
    .X(net433));
 sky130_fd_sc_hd__a31o_1 c683 (.A1(net315),
    .A2(net29),
    .A3(net139),
    .B1(net842),
    .X(net434));
 sky130_fd_sc_hd__a31o_1 c684 (.A1(net243),
    .A2(net626),
    .A3(net215),
    .B1(net346),
    .X(net435));
 sky130_fd_sc_hd__a31o_1 c685 (.A1(net212),
    .A2(net315),
    .A3(net851),
    .B1(net829),
    .X(net436));
 sky130_fd_sc_hd__a41o_1 c686 (.A1(net137),
    .A2(net215),
    .A3(net724),
    .A4(net225),
    .B1(net571),
    .X(net437));
 sky130_fd_sc_hd__a41o_1 c687 (.A1(net124),
    .A2(net411),
    .A3(net816),
    .A4(net346),
    .B1(net123),
    .X(net438));
 sky130_fd_sc_hd__a31o_1 c688 (.A1(net322),
    .A2(net434),
    .A3(net562),
    .B1(net842),
    .X(net439));
 sky130_fd_sc_hd__a31o_1 c689 (.A1(net435),
    .A2(net343),
    .A3(net242),
    .B1(net829),
    .X(net440));
 sky130_fd_sc_hd__a21bo_1 c690 (.A1(net434),
    .A2(net317),
    .B1_N(net549),
    .X(net441));
 sky130_fd_sc_hd__mux4_1 c691 (.A0(net225),
    .A1(net412),
    .A2(net849),
    .A3(net543),
    .S0(net843),
    .S1(net609),
    .X(net442));
 sky130_fd_sc_hd__a31o_1 c692 (.A1(net308),
    .A2(net427),
    .A3(net656),
    .B1(net660),
    .X(net443));
 sky130_fd_sc_hd__a31o_1 c693 (.A1(net441),
    .A2(net211),
    .A3(net426),
    .B1(net829),
    .X(net444));
 sky130_fd_sc_hd__a31o_1 c694 (.A1(net423),
    .A2(net902),
    .A3(net142),
    .B1(net562),
    .X(net445));
 sky130_fd_sc_hd__a21bo_1 c695 (.A1(net311),
    .A2(net807),
    .B1_N(net902),
    .X(net446));
 sky130_fd_sc_hd__a31o_1 c696 (.A1(net434),
    .A2(net823),
    .A3(net342),
    .B1(net435),
    .X(net447));
 sky130_fd_sc_hd__mux4_1 c697 (.A0(net442),
    .A1(net334),
    .A2(net412),
    .A3(net227),
    .S0(net212),
    .S1(net549),
    .X(net448));
 sky130_fd_sc_hd__a31o_1 c698 (.A1(net902),
    .A2(net437),
    .A3(net311),
    .B1(net571),
    .X(net449));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(net446),
    .A1(net139),
    .A2(net441),
    .A3(net571),
    .S0(net607),
    .S1(net609),
    .X(net450));
 sky130_fd_sc_hd__a31o_2 c700 (.A1(net427),
    .A2(net139),
    .A3(net548),
    .B1(net571),
    .X(net451));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(net444),
    .A1(net660),
    .A2(net817),
    .A3(net426),
    .S0(net142),
    .S1(net609),
    .X(net452));
 sky130_fd_sc_hd__a31o_1 c702 (.A1(net215),
    .A2(net883),
    .A3(net438),
    .B1(net543),
    .X(net453));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(net443),
    .A1(net453),
    .A2(net436),
    .A3(net415),
    .S0(net243),
    .S1(net608),
    .X(net454));
 sky130_fd_sc_hd__a41o_1 c704 (.A1(net310),
    .A2(net835),
    .A3(net723),
    .A4(net249),
    .B1(net817),
    .X(net455));
 sky130_fd_sc_hd__sdfbbn_1 c705 (.CLK_N(clknet_2_0__leaf_clk),
    .D(net416),
    .RESET_B(net660),
    .SCD(net453),
    .SCE(net847),
    .SET_B(net893),
    .Q(net457),
    .Q_N(net456));
 sky130_fd_sc_hd__mux4_1 c706 (.A0(net242),
    .A1(net142),
    .A2(net311),
    .A3(net724),
    .S0(net368),
    .S1(net622),
    .X(net458));
 sky130_fd_sc_hd__mux4_1 c707 (.A0(net671),
    .A1(net314),
    .A2(net265),
    .A3(net227),
    .S0(net723),
    .S1(net805),
    .X(net459));
 sky130_fd_sc_hd__mux4_2 c708 (.A0(net148),
    .A1(net123),
    .A2(net456),
    .A3(net817),
    .S0(net841),
    .S1(net622),
    .X(net460));
 sky130_fd_sc_hd__a41o_1 c709 (.A1(net891),
    .A2(net458),
    .A3(net415),
    .A4(net346),
    .B1(net544),
    .X(net461));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net438),
    .A1(net249),
    .A2(net451),
    .A3(net415),
    .S0(net882),
    .S1(net607),
    .X(net462));
 sky130_fd_sc_hd__mux4_2 c711 (.A0(net228),
    .A1(net131),
    .A2(net436),
    .A3(net850),
    .S0(net346),
    .S1(net626),
    .X(net463));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net807),
    .A1(net334),
    .A2(net872),
    .A3(net805),
    .S0(net848),
    .S1(net841),
    .X(net464));
 sky130_fd_sc_hd__a41o_1 c713 (.A1(net368),
    .A2(net428),
    .A3(net148),
    .A4(net548),
    .B1(net611),
    .X(net465));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(net465),
    .A1(net410),
    .A2(net807),
    .A3(net884),
    .S0(net314),
    .S1(net412),
    .X(net466));
 sky130_fd_sc_hd__a41o_1 c715 (.A1(net357),
    .A2(net123),
    .A3(net429),
    .A4(net416),
    .B1(clknet_1_0__leaf_net367),
    .X(net467));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(clknet_1_0__leaf_net367),
    .A1(net429),
    .A2(net671),
    .A3(net660),
    .S0(net850),
    .S1(clknet_1_0__leaf_net614),
    .X(net468));
 sky130_fd_sc_hd__a41o_1 c717 (.A1(net222),
    .A2(net460),
    .A3(net428),
    .A4(net726),
    .B1(clknet_1_0__leaf_net615),
    .X(net469));
 sky130_fd_sc_hd__sdfbbn_1 c718 (.CLK_N(clknet_2_0__leaf_clk),
    .D(net334),
    .RESET_B(net824),
    .SCD(clknet_1_0__leaf_net162),
    .SCE(net457),
    .SET_B(net829),
    .Q(net471),
    .Q_N(net470));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net225),
    .A1(net469),
    .A2(net444),
    .A3(net470),
    .S0(net851),
    .S1(net656),
    .X(net472));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net346),
    .A1(net891),
    .A2(net465),
    .A3(net819),
    .S0(net851),
    .S1(clknet_1_0__leaf_net614),
    .X(net473));
 sky130_fd_sc_hd__a41o_1 c721 (.A1(net462),
    .A2(net471),
    .A3(net660),
    .A4(net671),
    .B1(clknet_1_0__leaf_net614),
    .X(net474));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net412),
    .A1(net470),
    .A2(net222),
    .A3(net880),
    .S0(net743),
    .S1(clknet_1_0__leaf_net615),
    .X(net475));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net453),
    .A1(net227),
    .A2(net460),
    .A3(net415),
    .S0(net317),
    .S1(net433),
    .X(net476));
 sky130_fd_sc_hd__a41o_1 c724 (.A1(net437),
    .A2(net452),
    .A3(net886),
    .A4(clknet_1_0__leaf_net473),
    .B1(clknet_1_0__leaf_net614),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net436),
    .A1(net471),
    .A2(net410),
    .A3(net605),
    .S0(net611),
    .S1(clknet_1_1__leaf_net614),
    .X(net729));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net318),
    .A1(net439),
    .A2(net848),
    .A3(net353),
    .S0(net451),
    .S1(net842),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(clknet_1_0__leaf_net473),
    .A1(net37),
    .A2(net847),
    .A3(clknet_1_0__leaf_net162),
    .S0(net456),
    .S1(clknet_1_0__leaf_net615),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net455),
    .A1(net450),
    .A2(net806),
    .A3(net835),
    .S0(net609),
    .S1(net622),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(net859),
    .A1(clknet_1_1__leaf_net475),
    .A2(net731),
    .A3(net835),
    .S0(net702),
    .S1(net759),
    .X(net481));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net410),
    .A1(net738),
    .A2(net884),
    .A3(net605),
    .S0(net609),
    .S1(net759),
    .X(net482));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net354),
    .A1(net173),
    .A2(net629),
    .A3(net544),
    .S0(net619),
    .S1(net622),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(net878),
    .A1(net457),
    .A2(net59),
    .A3(net683),
    .S0(net667),
    .S1(net616),
    .X(net484));
 sky130_fd_sc_hd__mux4_2 c733 (.A0(net668),
    .A1(net805),
    .A2(net68),
    .A3(net848),
    .S0(net822),
    .S1(net623),
    .X(net785));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(net484),
    .A1(net806),
    .A2(net641),
    .A3(net605),
    .S0(net618),
    .S1(net623),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net629),
    .A1(net40),
    .A2(net805),
    .A3(net738),
    .S0(net608),
    .S1(net623),
    .X(net486));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(net850),
    .A1(net466),
    .A2(net460),
    .A3(net723),
    .S0(net544),
    .S1(net623),
    .X(net487));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net307),
    .A1(net457),
    .A2(clknet_1_0__leaf_net370),
    .A3(net816),
    .S0(net702),
    .S1(net842),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net668),
    .A1(net71),
    .A2(net667),
    .A3(net142),
    .S0(net485),
    .S1(net815),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(net433),
    .A1(net59),
    .A2(net37),
    .A3(net439),
    .S0(net815),
    .S1(net460),
    .X(net490));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(net415),
    .A1(net353),
    .A2(net478),
    .A3(net850),
    .S0(net456),
    .S1(net623),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(net451),
    .A1(net486),
    .A2(net624),
    .A3(net71),
    .S0(net723),
    .S1(net606),
    .X(net492));
 sky130_fd_sc_hd__mux4_2 c742 (.A0(net129),
    .A1(net415),
    .A2(net410),
    .A3(net843),
    .S0(net607),
    .S1(net623),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(net491),
    .A1(clknet_1_0__leaf_net162),
    .A2(net692),
    .A3(net439),
    .S0(net785),
    .S1(net451),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(clknet_1_0__leaf_net475),
    .A1(net459),
    .A2(net173),
    .A3(clknet_1_1__leaf_net473),
    .S0(net40),
    .S1(net606),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(clknet_1_0__leaf_net162),
    .A1(net266),
    .A2(net463),
    .A3(net656),
    .S0(net611),
    .S1(net617),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net317),
    .A1(net701),
    .A2(net439),
    .A3(clknet_1_0__leaf_net615),
    .S0(net617),
    .S1(net623),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(net312),
    .A1(net497),
    .A2(net626),
    .A3(net616),
    .S0(net622),
    .S1(net623),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net373),
    .A1(net266),
    .A2(net393),
    .A3(net645),
    .S0(net641),
    .S1(net816),
    .X(net499));
 sky130_fd_sc_hd__mux4_2 c749 (.A0(net810),
    .A1(net406),
    .A2(net812),
    .A3(net629),
    .S0(net463),
    .S1(net613),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(net489),
    .A1(net293),
    .A2(net482),
    .A3(net681),
    .S0(net842),
    .S1(net608),
    .X(net501));
 sky130_fd_sc_hd__mux4_2 c751 (.A0(net37),
    .A1(net701),
    .A2(net498),
    .A3(net500),
    .S0(net835),
    .S1(net731),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net424),
    .A1(net354),
    .A2(net873),
    .A3(net886),
    .S0(net805),
    .S1(net842),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net84),
    .A1(net815),
    .A2(net493),
    .A3(net827),
    .S0(net844),
    .S1(net743),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net667),
    .A1(net681),
    .A2(net738),
    .A3(net600),
    .S0(net743),
    .S1(net617),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net624),
    .A1(net187),
    .A2(net668),
    .A3(net876),
    .S0(net744),
    .S1(net613),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net506),
    .A1(net830),
    .A2(net392),
    .A3(net629),
    .S0(net848),
    .S1(net611),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net819),
    .A1(net460),
    .A2(net480),
    .A3(net667),
    .S0(net194),
    .S1(net843),
    .X(net508));
 sky130_fd_sc_hd__mux4_2 c758 (.A0(net835),
    .A1(net40),
    .A2(net398),
    .A3(net173),
    .S0(net600),
    .S1(net822),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net722),
    .A1(net407),
    .A2(net641),
    .A3(net877),
    .S0(net597),
    .S1(net844),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net265),
    .A1(net187),
    .A2(net645),
    .A3(net600),
    .S0(net606),
    .S1(net611),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net343),
    .A1(clknet_1_1__leaf_net370),
    .A2(net835),
    .A3(net722),
    .S0(net724),
    .S1(net616),
    .X(net512));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net505),
    .A1(net656),
    .A2(net815),
    .A3(net609),
    .S0(net611),
    .S1(net613),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(clknet_1_0__leaf_net255),
    .A1(net194),
    .A2(net485),
    .A3(clknet_1_0__leaf_net512),
    .S0(net511),
    .S1(net744),
    .X(net514));
 sky130_fd_sc_hd__mux4_1 c764 (.A0(net692),
    .A1(net68),
    .A2(net108),
    .A3(net842),
    .S0(net759),
    .S1(clknet_1_1__leaf_net615),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c765 (.A0(net681),
    .A1(net624),
    .A2(net511),
    .A3(net738),
    .S0(clknet_1_1__leaf_net512),
    .S1(net600),
    .X(net516));
 sky130_fd_sc_hd__mux4_1 c766 (.A0(net702),
    .A1(clknet_1_0__leaf_net400),
    .A2(net492),
    .A3(net488),
    .S0(net597),
    .S1(net619),
    .X(net517));
 sky130_fd_sc_hd__mux4_1 c767 (.A0(net683),
    .A1(net698),
    .A2(net905),
    .A3(net515),
    .S0(net817),
    .S1(net609),
    .X(net518));
 sky130_fd_sc_hd__mux4_1 c768 (.A0(net513),
    .A1(net117),
    .A2(net667),
    .A3(net517),
    .S0(net657),
    .S1(net617),
    .X(net519));
 sky130_fd_sc_hd__mux4_1 c769 (.A0(net429),
    .A1(net519),
    .A2(net518),
    .A3(net625),
    .S0(clknet_1_1__leaf_net615),
    .S1(net619),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 merge790 (.A0(net169),
    .A1(clknet_1_1__leaf_net162),
    .A2(net694),
    .A3(net171),
    .S0(net755),
    .S1(net821),
    .X(net521));
 sky130_fd_sc_hd__a41o_1 merge791 (.A1(net244),
    .A2(clknet_1_0__leaf_net161),
    .A3(net625),
    .A4(net121),
    .B1(net246),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 merge792 (.A0(net55),
    .A1(net74),
    .A2(net810),
    .A3(net92),
    .S0(net86),
    .S1(net93),
    .X(net523));
 sky130_fd_sc_hd__mux4_1 merge793 (.A0(net320),
    .A1(net634),
    .A2(net330),
    .A3(net331),
    .S0(net847),
    .S1(net829),
    .X(net524));
 sky130_fd_sc_hd__mux4_2 merge794 (.A0(net258),
    .A1(net132),
    .A2(net761),
    .A3(net708),
    .S0(net93),
    .S1(net180),
    .X(net525));
 sky130_fd_sc_hd__mux4_1 merge795 (.A0(net330),
    .A1(net866),
    .A2(net311),
    .A3(net233),
    .S0(net232),
    .S1(net767),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 merge796 (.A0(net74),
    .A1(net77),
    .A2(net79),
    .A3(net88),
    .S0(net95),
    .S1(net698),
    .X(net527));
 sky130_fd_sc_hd__mux4_1 merge797 (.A0(clknet_1_1__leaf_net162),
    .A1(net47),
    .A2(net158),
    .A3(net155),
    .S0(net757),
    .S1(net169),
    .X(net528));
 sky130_fd_sc_hd__xnor2_1 merge798 (.A(net164),
    .B(net528),
    .Y(net529));
 sky130_fd_sc_hd__xnor2_1 merge799 (.A(net174),
    .B(net521),
    .Y(net530));
 sky130_fd_sc_hd__xnor2_1 merge800 (.A(net285),
    .B(net269),
    .Y(net531));
 sky130_fd_sc_hd__xnor2_1 merge801 (.A(net235),
    .B(net241),
    .Y(net532));
 sky130_fd_sc_hd__xnor2_1 merge802 (.A(net467),
    .B(net474),
    .Y(net533));
 sky130_fd_sc_hd__xnor2_1 merge803 (.A(net349),
    .B(net350),
    .Y(net534));
 sky130_fd_sc_hd__xnor2_1 merge804 (.A(net94),
    .B(net523),
    .Y(net535));
 sky130_fd_sc_hd__xnor2_1 merge805 (.A(net186),
    .B(net202),
    .Y(net536));
 sky130_fd_sc_hd__xnor2_1 merge806 (.A(net391),
    .B(net396),
    .Y(net537));
 sky130_fd_sc_hd__xnor2_1 merge807 (.A(net287),
    .B(net294),
    .Y(net538));
 sky130_fd_sc_hd__xnor2_1 merge808 (.A(net102),
    .B(net104),
    .Y(net539));
 sky130_fd_sc_hd__xnor2_1 merge809 (.A(net481),
    .B(net487),
    .Y(net540));
 sky130_fd_sc_hd__xnor2_1 merge810 (.A(net520),
    .B(net499),
    .Y(net541));
 sky130_fd_sc_hd__xnor2_1 merge811 (.A(net376),
    .B(net379),
    .Y(net542));
 sky130_fd_sc_hd__dfrbp_2 merge812 (.CLK(clknet_2_0__leaf_clk),
    .D(net425),
    .RESET_B(net430),
    .Q(net544),
    .Q_N(net543));
 sky130_fd_sc_hd__xnor2_1 merge813 (.A(net345),
    .B(net332),
    .Y(net545));
 sky130_fd_sc_hd__xnor2_1 merge814 (.A(net253),
    .B(net256),
    .Y(net546));
 sky130_fd_sc_hd__xnor2_1 merge815 (.A(net75),
    .B(net527),
    .Y(net547));
 sky130_fd_sc_hd__dfrbp_1 merge816 (.CLK(clknet_2_0__leaf_clk),
    .D(net440),
    .RESET_B(net447),
    .Q(net549),
    .Q_N(net548));
 sky130_fd_sc_hd__xnor2_1 merge817 (.A(net264),
    .B(net522),
    .Y(net550));
 sky130_fd_sc_hd__xnor2_1 merge818 (.A(net157),
    .B(net163),
    .Y(net551));
 sky130_fd_sc_hd__xnor2_1 merge819 (.A(net401),
    .B(net409),
    .Y(net552));
 sky130_fd_sc_hd__xnor2_1 merge820 (.A(net541),
    .B(net516),
    .Y(net553));
 sky130_fd_sc_hd__xnor2_1 merge821 (.A(net101),
    .B(net103),
    .Y(net554));
 sky130_fd_sc_hd__xnor2_1 merge822 (.A(net380),
    .B(net306),
    .Y(net555));
 sky130_fd_sc_hd__xnor2_1 merge823 (.A(net361),
    .B(net389),
    .Y(net556));
 sky130_fd_sc_hd__xnor2_1 merge824 (.A(net304),
    .B(net404),
    .Y(net557));
 sky130_fd_sc_hd__xnor2_1 merge825 (.A(net364),
    .B(net525),
    .Y(net558));
 sky130_fd_sc_hd__xnor2_1 merge826 (.A(net76),
    .B(net78),
    .Y(net559));
 sky130_fd_sc_hd__xnor2_1 merge827 (.A(net539),
    .B(net96),
    .Y(net560));
 sky130_fd_sc_hd__xnor2_1 merge828 (.A(net288),
    .B(net297),
    .Y(net561));
 sky130_fd_sc_hd__dfrtn_1 merge829 (.CLK_N(clknet_2_0__leaf_clk),
    .D(net347),
    .RESET_B(net524),
    .Q(net562));
 sky130_fd_sc_hd__xnor2_1 merge830 (.A(net494),
    .B(net514),
    .Y(net563));
 sky130_fd_sc_hd__xnor2_1 merge831 (.A(net495),
    .B(net510),
    .Y(net564));
 sky130_fd_sc_hd__xnor2_2 merge832 (.A(net501),
    .B(net502),
    .Y(net565));
 sky130_fd_sc_hd__xnor2_1 merge833 (.A(net564),
    .B(net286),
    .Y(net566));
 sky130_fd_sc_hd__xnor2_1 merge834 (.A(net83),
    .B(net529),
    .Y(net567));
 sky130_fd_sc_hd__xnor2_1 merge835 (.A(net82),
    .B(net547),
    .Y(net568));
 sky130_fd_sc_hd__dfrtp_1 merge836 (.CLK(clknet_2_2__leaf_clk),
    .D(net526),
    .RESET_B(net352),
    .Q(net569));
 sky130_fd_sc_hd__xnor2_2 merge837 (.A(net509),
    .B(net504),
    .Y(net570));
 sky130_fd_sc_hd__dfrtp_2 merge838 (.CLK(clknet_2_0__leaf_clk),
    .D(net448),
    .RESET_B(net431),
    .Q(net571));
 sky130_fd_sc_hd__dfrtp_2 merge839 (.CLK(clknet_2_2__leaf_clk),
    .D(net559),
    .RESET_B(net567),
    .Q(net572));
 sky130_fd_sc_hd__dfsbp_1 merge840 (.CLK(clknet_2_0__leaf_clk),
    .D(net344),
    .SET_B(net545),
    .Q(net574),
    .Q_N(net573));
 sky130_fd_sc_hd__xnor2_1 merge841 (.A(net280),
    .B(net283),
    .Y(net575));
 sky130_fd_sc_hd__xnor2_1 merge842 (.A(net531),
    .B(net546),
    .Y(net576));
 sky130_fd_sc_hd__xnor2_1 merge843 (.A(net535),
    .B(net554),
    .Y(net577));
 sky130_fd_sc_hd__xnor2_1 merge844 (.A(net461),
    .B(net477),
    .Y(net578));
 sky130_fd_sc_hd__xnor2_1 merge845 (.A(net508),
    .B(net302),
    .Y(net579));
 sky130_fd_sc_hd__xnor2_1 merge846 (.A(net303),
    .B(net538),
    .Y(net580));
 sky130_fd_sc_hd__xnor2_1 merge847 (.A(net472),
    .B(net563),
    .Y(net581));
 sky130_fd_sc_hd__xnor2_1 merge848 (.A(net184),
    .B(net530),
    .Y(net582));
 sky130_fd_sc_hd__xnor2_1 merge849 (.A(net536),
    .B(net160),
    .Y(net583));
 sky130_fd_sc_hd__xnor2_1 merge850 (.A(net557),
    .B(net291),
    .Y(net584));
 sky130_fd_sc_hd__xnor2_1 merge851 (.A(net377),
    .B(net552),
    .Y(net585));
 sky130_fd_sc_hd__xnor2_1 merge852 (.A(net468),
    .B(net405),
    .Y(net586));
 sky130_fd_sc_hd__xnor2_1 merge853 (.A(net540),
    .B(net496),
    .Y(net587));
 sky130_fd_sc_hd__xnor2_1 merge854 (.A(net555),
    .B(net542),
    .Y(net588));
 sky130_fd_sc_hd__xnor2_1 merge855 (.A(net386),
    .B(net537),
    .Y(net589));
 sky130_fd_sc_hd__xnor2_2 merge856 (.A(net402),
    .B(net570),
    .Y(net590));
 sky130_fd_sc_hd__xnor2_1 merge857 (.A(net355),
    .B(net533),
    .Y(net591));
 sky130_fd_sc_hd__dfsbp_1 merge858 (.CLK(clknet_2_3__leaf_clk),
    .D(net397),
    .SET_B(net284),
    .Q(net593),
    .Q_N(net592));
 sky130_fd_sc_hd__xnor2_1 merge859 (.A(net565),
    .B(net534),
    .Y(net594));
 sky130_fd_sc_hd__xnor2_1 merge860 (.A(net476),
    .B(net556),
    .Y(net595));
 sky130_fd_sc_hd__xnor2_1 merge861 (.A(net479),
    .B(net553),
    .Y(net596));
 sky130_fd_sc_hd__dfstp_2 merge862 (.CLK(clknet_2_1__leaf_clk),
    .D(net362),
    .SET_B(net507),
    .Q(net597));
 sky130_fd_sc_hd__xnor2_1 merge863 (.A(net550),
    .B(net575),
    .Y(net598));
 sky130_fd_sc_hd__xnor2_1 merge864 (.A(net560),
    .B(net551),
    .Y(net599));
 sky130_fd_sc_hd__dfstp_2 merge865 (.CLK(clknet_2_1__leaf_clk),
    .D(net579),
    .SET_B(net503),
    .Q(net600));
 sky130_fd_sc_hd__dfstp_1 merge866 (.CLK(clknet_2_2__leaf_clk),
    .D(net582),
    .SET_B(net568),
    .Q(net601));
 sky130_fd_sc_hd__dlrbn_1 merge867 (.D(net598),
    .GATE_N(clknet_2_2__leaf_clk),
    .RESET_B(net532),
    .Q(net753),
    .Q_N(net602));
 sky130_fd_sc_hd__dlrbn_2 merge868 (.D(net576),
    .GATE_N(clknet_2_2__leaf_clk),
    .RESET_B(net181),
    .Q(net603),
    .Q_N(net734));
 sky130_fd_sc_hd__dlrbp_1 merge869 (.D(net369),
    .GATE(clknet_2_2__leaf_clk),
    .RESET_B(net558),
    .Q(net605),
    .Q_N(net604));
 sky130_fd_sc_hd__dlrbp_1 merge870 (.D(net445),
    .GATE(clknet_2_1__leaf_clk),
    .RESET_B(net490),
    .Q(net607),
    .Q_N(net606));
 sky130_fd_sc_hd__dlrtn_4 merge871 (.D(net449),
    .GATE_N(clknet_2_3__leaf_clk),
    .RESET_B(net589),
    .Q(net608));
 sky130_fd_sc_hd__dlrtn_4 merge872 (.D(net432),
    .GATE_N(clknet_2_1__leaf_clk),
    .RESET_B(net596),
    .Q(net609));
 sky130_fd_sc_hd__dlrtn_4 merge873 (.D(net585),
    .GATE_N(clknet_2_3__leaf_clk),
    .RESET_B(net588),
    .Q(net759));
 sky130_fd_sc_hd__xnor2_1 merge874 (.A(net561),
    .B(net365),
    .Y(net610));
 sky130_fd_sc_hd__dlrtp_4 merge875 (.GATE(clknet_2_2__leaf_clk),
    .RESET_B(net165),
    .Q(net748));
 sky130_fd_sc_hd__dlrtp_4 merge876 (.D(net591),
    .GATE(clknet_2_0__leaf_clk),
    .RESET_B(net594),
    .Q(net743));
 sky130_fd_sc_hd__dlrtp_4 merge877 (.D(net578),
    .GATE(clknet_2_1__leaf_clk),
    .RESET_B(net590),
    .Q(net611));
 sky130_fd_sc_hd__edfxbp_1 merge878 (.CLK(clknet_2_3__leaf_clk),
    .D(net580),
    .DE(net584),
    .Q(net613),
    .Q_N(net612));
 sky130_fd_sc_hd__edfxtp_1 merge879 (.CLK(clknet_2_3__leaf_clk),
    .D(net577),
    .DE(net610),
    .Q(net801));
 sky130_fd_sc_hd__sdlclkp_1 merge880 (.CLK(clknet_2_1__leaf_clk),
    .GATE(net464),
    .SCE(net595),
    .GCLK(net614));
 sky130_fd_sc_hd__sdlclkp_2 merge881 (.CLK(clknet_2_2__leaf_clk),
    .GATE(net583),
    .SCE(net599),
    .GCLK(net799));
 sky130_fd_sc_hd__sdlclkp_4 merge882 (.CLK(clknet_2_1__leaf_clk),
    .GATE(net586),
    .SCE(net581),
    .GCLK(net615));
 sky130_fd_sc_hd__dfrbp_2 merge883 (.CLK(clknet_2_1__leaf_clk),
    .D(net587),
    .RESET_B(net566),
    .Q(net617),
    .Q_N(net616));
 sky130_fd_sc_hd__dfxbp_1 s884 (.CLK(clknet_2_2__leaf_clk),
    .D(net363),
    .Q(net619),
    .Q_N(net618));
 sky130_fd_sc_hd__dfxbp_1 s885 (.CLK(clknet_2_3__leaf_clk),
    .D(net399),
    .Q(net621),
    .Q_N(net620));
 sky130_fd_sc_hd__dfxtp_2 s886 (.CLK(clknet_2_0__leaf_clk),
    .D(net454),
    .Q(net622));
 sky130_fd_sc_hd__dfxtp_2 s887 (.CLK(clknet_2_1__leaf_clk),
    .D(net483),
    .Q(net623));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_6 input1 (.A(in0),
    .X(net182));
 sky130_fd_sc_hd__buf_2 input2 (.A(in1),
    .X(net624));
 sky130_fd_sc_hd__buf_6 input3 (.A(in10),
    .X(net625));
 sky130_fd_sc_hd__buf_4 input4 (.A(in11),
    .X(net626));
 sky130_fd_sc_hd__buf_1 input5 (.A(in12),
    .X(net627));
 sky130_fd_sc_hd__buf_4 input6 (.A(in13),
    .X(net628));
 sky130_fd_sc_hd__buf_4 input7 (.A(in14),
    .X(net629));
 sky130_fd_sc_hd__buf_2 input8 (.A(in15),
    .X(net630));
 sky130_fd_sc_hd__buf_4 input9 (.A(in16),
    .X(net631));
 sky130_fd_sc_hd__buf_2 input10 (.A(in17),
    .X(net632));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(in18),
    .X(net633));
 sky130_fd_sc_hd__buf_4 input12 (.A(in19),
    .X(net634));
 sky130_fd_sc_hd__clkbuf_8 input13 (.A(in2),
    .X(net635));
 sky130_fd_sc_hd__buf_4 input14 (.A(in20),
    .X(net636));
 sky130_fd_sc_hd__buf_4 input15 (.A(in21),
    .X(net637));
 sky130_fd_sc_hd__buf_2 input16 (.A(in22),
    .X(net638));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(in23),
    .X(net639));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(in24),
    .X(net640));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(in25),
    .X(net641));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(in26),
    .X(net642));
 sky130_fd_sc_hd__buf_2 input21 (.A(in27),
    .X(net643));
 sky130_fd_sc_hd__dlymetal6s2s_1 input22 (.A(in28),
    .X(net644));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(in29),
    .X(net645));
 sky130_fd_sc_hd__buf_4 input24 (.A(in3),
    .X(net646));
 sky130_fd_sc_hd__buf_2 input25 (.A(in30),
    .X(net647));
 sky130_fd_sc_hd__buf_2 input26 (.A(in31),
    .X(net648));
 sky130_fd_sc_hd__buf_2 input27 (.A(in32),
    .X(net649));
 sky130_fd_sc_hd__buf_4 input28 (.A(in33),
    .X(net650));
 sky130_fd_sc_hd__buf_4 input29 (.A(in34),
    .X(net651));
 sky130_fd_sc_hd__dlymetal6s2s_1 input30 (.A(in35),
    .X(net652));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(in36),
    .X(net653));
 sky130_fd_sc_hd__buf_2 input32 (.A(in37),
    .X(net654));
 sky130_fd_sc_hd__dlymetal6s2s_1 input33 (.A(in38),
    .X(net655));
 sky130_fd_sc_hd__buf_4 input34 (.A(in39),
    .X(net656));
 sky130_fd_sc_hd__buf_8 input35 (.A(in4),
    .X(net657));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(in40),
    .X(net658));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(in41),
    .X(net659));
 sky130_fd_sc_hd__clkbuf_4 input38 (.A(in42),
    .X(net660));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(in43),
    .X(net661));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(in44),
    .X(net662));
 sky130_fd_sc_hd__buf_1 input41 (.A(in45),
    .X(net663));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(in46),
    .X(net664));
 sky130_fd_sc_hd__buf_2 input43 (.A(in47),
    .X(net665));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(in48),
    .X(net666));
 sky130_fd_sc_hd__buf_4 input45 (.A(in49),
    .X(net667));
 sky130_fd_sc_hd__clkbuf_8 input46 (.A(in5),
    .X(net668));
 sky130_fd_sc_hd__buf_1 input47 (.A(in50),
    .X(net669));
 sky130_fd_sc_hd__buf_1 input48 (.A(in51),
    .X(net670));
 sky130_fd_sc_hd__buf_2 input49 (.A(in52),
    .X(net671));
 sky130_fd_sc_hd__clkbuf_4 input50 (.A(in53),
    .X(net672));
 sky130_fd_sc_hd__buf_2 input51 (.A(in54),
    .X(net673));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(in55),
    .X(net674));
 sky130_fd_sc_hd__buf_1 input53 (.A(in56),
    .X(net675));
 sky130_fd_sc_hd__buf_1 input54 (.A(in57),
    .X(net676));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(in58),
    .X(net677));
 sky130_fd_sc_hd__dlymetal6s2s_1 input56 (.A(in59),
    .X(net678));
 sky130_fd_sc_hd__clkbuf_8 input57 (.A(in6),
    .X(net679));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(in60),
    .X(net680));
 sky130_fd_sc_hd__clkbuf_4 input59 (.A(in61),
    .X(net681));
 sky130_fd_sc_hd__dlymetal6s2s_1 input60 (.A(in62),
    .X(net682));
 sky130_fd_sc_hd__buf_4 input61 (.A(in63),
    .X(net683));
 sky130_fd_sc_hd__dlymetal6s2s_1 input62 (.A(in64),
    .X(net684));
 sky130_fd_sc_hd__buf_4 input63 (.A(in65),
    .X(net685));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(in66),
    .X(net686));
 sky130_fd_sc_hd__buf_1 input65 (.A(in67),
    .X(net687));
 sky130_fd_sc_hd__buf_1 input66 (.A(in68),
    .X(net688));
 sky130_fd_sc_hd__buf_1 input67 (.A(in69),
    .X(net689));
 sky130_fd_sc_hd__buf_4 input68 (.A(in7),
    .X(net690));
 sky130_fd_sc_hd__buf_2 input69 (.A(in70),
    .X(net691));
 sky130_fd_sc_hd__buf_2 input70 (.A(in71),
    .X(net692));
 sky130_fd_sc_hd__clkbuf_2 input71 (.A(in72),
    .X(net693));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(in73),
    .X(net694));
 sky130_fd_sc_hd__buf_1 input73 (.A(in74),
    .X(net695));
 sky130_fd_sc_hd__clkbuf_2 input74 (.A(in75),
    .X(net696));
 sky130_fd_sc_hd__buf_2 input75 (.A(in76),
    .X(net697));
 sky130_fd_sc_hd__clkbuf_4 input76 (.A(in77),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_4 input77 (.A(in78),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_2 input78 (.A(in79),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(in8),
    .X(net701));
 sky130_fd_sc_hd__buf_4 input80 (.A(in80),
    .X(net702));
 sky130_fd_sc_hd__clkbuf_2 input81 (.A(in81),
    .X(net703));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(in82),
    .X(net704));
 sky130_fd_sc_hd__buf_1 input83 (.A(in83),
    .X(net705));
 sky130_fd_sc_hd__clkbuf_2 input84 (.A(in84),
    .X(net706));
 sky130_fd_sc_hd__dlymetal6s2s_1 input85 (.A(in85),
    .X(net707));
 sky130_fd_sc_hd__dlymetal6s2s_1 input86 (.A(in86),
    .X(net708));
 sky130_fd_sc_hd__buf_2 input87 (.A(in87),
    .X(net709));
 sky130_fd_sc_hd__dlymetal6s2s_1 input88 (.A(in88),
    .X(net710));
 sky130_fd_sc_hd__buf_1 input89 (.A(in89),
    .X(net711));
 sky130_fd_sc_hd__buf_4 input90 (.A(in9),
    .X(net712));
 sky130_fd_sc_hd__clkbuf_4 input91 (.A(in90),
    .X(net713));
 sky130_fd_sc_hd__buf_1 input92 (.A(in91),
    .X(net714));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(in92),
    .X(net715));
 sky130_fd_sc_hd__dlymetal6s2s_1 input94 (.A(in93),
    .X(net716));
 sky130_fd_sc_hd__clkbuf_2 input95 (.A(in94),
    .X(net717));
 sky130_fd_sc_hd__buf_1 input96 (.A(in95),
    .X(net718));
 sky130_fd_sc_hd__dlymetal6s2s_1 input97 (.A(in96),
    .X(net719));
 sky130_fd_sc_hd__buf_1 input98 (.A(in97),
    .X(net720));
 sky130_fd_sc_hd__clkbuf_2 input99 (.A(in98),
    .X(net721));
 sky130_fd_sc_hd__clkbuf_4 input100 (.A(in99),
    .X(net722));
 sky130_fd_sc_hd__buf_2 output101 (.A(net723),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output102 (.A(net724),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output103 (.A(net817),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output104 (.A(net726),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output105 (.A(net806),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output106 (.A(net876),
    .X(out14));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(net729),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output108 (.A(net868),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output109 (.A(net731),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output110 (.A(net885),
    .X(out19));
 sky130_fd_sc_hd__clkbuf_4 output111 (.A(net733),
    .X(out2));
 sky130_fd_sc_hd__clkbuf_4 output112 (.A(net734),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output113 (.A(net735),
    .X(out21));
 sky130_fd_sc_hd__clkbuf_4 output114 (.A(net736),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output115 (.A(net737),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output116 (.A(net738),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output117 (.A(net739),
    .X(out25));
 sky130_fd_sc_hd__buf_2 output118 (.A(net886),
    .X(out27));
 sky130_fd_sc_hd__clkbuf_1 output119 (.A(net741),
    .X(out28));
 sky130_fd_sc_hd__clkbuf_1 output120 (.A(clknet_1_1__leaf_net742),
    .X(out29));
 sky130_fd_sc_hd__buf_2 output121 (.A(net743),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output122 (.A(net823),
    .X(out30));
 sky130_fd_sc_hd__clkbuf_4 output123 (.A(net745),
    .X(out31));
 sky130_fd_sc_hd__clkbuf_4 output124 (.A(net746),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output125 (.A(net747),
    .X(out36));
 sky130_fd_sc_hd__buf_2 output126 (.A(net822),
    .X(out37));
 sky130_fd_sc_hd__buf_2 output127 (.A(net749),
    .X(out38));
 sky130_fd_sc_hd__clkbuf_4 output128 (.A(net750),
    .X(out39));
 sky130_fd_sc_hd__buf_2 output129 (.A(net751),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output130 (.A(net752),
    .X(out41));
 sky130_fd_sc_hd__buf_2 output131 (.A(net843),
    .X(out42));
 sky130_fd_sc_hd__clkbuf_4 output132 (.A(net754),
    .X(out44));
 sky130_fd_sc_hd__clkbuf_4 output133 (.A(net755),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output134 (.A(net756),
    .X(out46));
 sky130_fd_sc_hd__clkbuf_4 output135 (.A(net757),
    .X(out48));
 sky130_fd_sc_hd__clkbuf_4 output136 (.A(net758),
    .X(out49));
 sky130_fd_sc_hd__buf_2 output137 (.A(net759),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output138 (.A(net760),
    .X(out51));
 sky130_fd_sc_hd__buf_2 output139 (.A(net761),
    .X(out52));
 sky130_fd_sc_hd__clkbuf_4 output140 (.A(net762),
    .X(out53));
 sky130_fd_sc_hd__clkbuf_4 output141 (.A(net763),
    .X(out54));
 sky130_fd_sc_hd__clkbuf_4 output142 (.A(net764),
    .X(out55));
 sky130_fd_sc_hd__clkbuf_4 output143 (.A(net765),
    .X(out57));
 sky130_fd_sc_hd__clkbuf_1 output144 (.A(clknet_1_1__leaf_net766),
    .X(out58));
 sky130_fd_sc_hd__buf_2 output145 (.A(net767),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output146 (.A(net768),
    .X(out60));
 sky130_fd_sc_hd__clkbuf_1 output147 (.A(clknet_1_1__leaf_net769),
    .X(out61));
 sky130_fd_sc_hd__clkbuf_4 output148 (.A(net770),
    .X(out62));
 sky130_fd_sc_hd__clkbuf_4 output149 (.A(net854),
    .X(out64));
 sky130_fd_sc_hd__clkbuf_4 output150 (.A(net772),
    .X(out65));
 sky130_fd_sc_hd__clkbuf_4 output151 (.A(net773),
    .X(out66));
 sky130_fd_sc_hd__clkbuf_4 output152 (.A(net774),
    .X(out67));
 sky130_fd_sc_hd__clkbuf_4 output153 (.A(net775),
    .X(out69));
 sky130_fd_sc_hd__clkbuf_4 output154 (.A(net776),
    .X(out70));
 sky130_fd_sc_hd__buf_2 output155 (.A(net777),
    .X(out71));
 sky130_fd_sc_hd__clkbuf_4 output156 (.A(net778),
    .X(out72));
 sky130_fd_sc_hd__clkbuf_4 output157 (.A(net779),
    .X(out73));
 sky130_fd_sc_hd__buf_2 output158 (.A(net780),
    .X(out75));
 sky130_fd_sc_hd__clkbuf_4 output159 (.A(net781),
    .X(out76));
 sky130_fd_sc_hd__clkbuf_4 output160 (.A(net782),
    .X(out77));
 sky130_fd_sc_hd__clkbuf_4 output161 (.A(net783),
    .X(out78));
 sky130_fd_sc_hd__clkbuf_4 output162 (.A(net784),
    .X(out79));
 sky130_fd_sc_hd__buf_2 output163 (.A(net785),
    .X(out8));
 sky130_fd_sc_hd__clkbuf_1 output164 (.A(clknet_1_1__leaf_net786),
    .X(out83));
 sky130_fd_sc_hd__buf_2 output165 (.A(net787),
    .X(out84));
 sky130_fd_sc_hd__clkbuf_4 output166 (.A(net788),
    .X(out85));
 sky130_fd_sc_hd__buf_2 output167 (.A(net789),
    .X(out86));
 sky130_fd_sc_hd__clkbuf_4 output168 (.A(net790),
    .X(out87));
 sky130_fd_sc_hd__clkbuf_4 output169 (.A(net840),
    .X(out88));
 sky130_fd_sc_hd__clkbuf_4 output170 (.A(net792),
    .X(out89));
 sky130_fd_sc_hd__clkbuf_1 output171 (.A(clknet_1_1__leaf_net793),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_4 output172 (.A(net794),
    .X(out90));
 sky130_fd_sc_hd__clkbuf_4 output173 (.A(net795),
    .X(out91));
 sky130_fd_sc_hd__buf_2 output174 (.A(net796),
    .X(out92));
 sky130_fd_sc_hd__buf_2 output175 (.A(net797),
    .X(out93));
 sky130_fd_sc_hd__buf_2 output176 (.A(net798),
    .X(out94));
 sky130_fd_sc_hd__clkbuf_1 output177 (.A(clknet_1_1__leaf_net799),
    .X(out95));
 sky130_fd_sc_hd__clkbuf_1 output178 (.A(clknet_1_0__leaf_net800),
    .X(out96));
 sky130_fd_sc_hd__clkbuf_4 output179 (.A(net801),
    .X(out97));
 sky130_fd_sc_hd__buf_2 output180 (.A(net802),
    .X(out98));
 sky130_fd_sc_hd__clkbuf_4 output181 (.A(net867),
    .X(out99));
 sky130_fd_sc_hd__buf_4 fanout182 (.A(net735),
    .X(net804));
 sky130_fd_sc_hd__buf_4 fanout183 (.A(net806),
    .X(net805));
 sky130_fd_sc_hd__clkbuf_4 fanout184 (.A(net727),
    .X(net806));
 sky130_fd_sc_hd__buf_4 fanout185 (.A(net216),
    .X(net807));
 sky130_fd_sc_hd__buf_4 fanout186 (.A(net733),
    .X(net808));
 sky130_fd_sc_hd__buf_4 fanout187 (.A(net203),
    .X(net809));
 sky130_fd_sc_hd__buf_4 fanout188 (.A(net69),
    .X(net810));
 sky130_fd_sc_hd__clkbuf_4 fanout189 (.A(net812),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_4 fanout190 (.A(net89),
    .X(net812));
 sky130_fd_sc_hd__buf_12 fanout191 (.A(net732),
    .X(net813));
 sky130_fd_sc_hd__buf_4 fanout192 (.A(net763),
    .X(net814));
 sky130_fd_sc_hd__buf_4 max_cap193 (.A(net110),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_8 fanout194 (.A(net117),
    .X(net816));
 sky130_fd_sc_hd__clkbuf_8 fanout195 (.A(net725),
    .X(net817));
 sky130_fd_sc_hd__buf_12 fanout196 (.A(net740),
    .X(net818));
 sky130_fd_sc_hd__buf_8 fanout197 (.A(net108),
    .X(net819));
 sky130_fd_sc_hd__buf_6 max_cap198 (.A(net27),
    .X(net820));
 sky130_fd_sc_hd__clkbuf_4 fanout199 (.A(net822),
    .X(net821));
 sky130_fd_sc_hd__buf_4 fanout200 (.A(net748),
    .X(net822));
 sky130_fd_sc_hd__buf_4 max_cap201 (.A(net744),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_8 fanout202 (.A(net107),
    .X(net824));
 sky130_fd_sc_hd__buf_12 fanout203 (.A(net827),
    .X(net825));
 sky130_fd_sc_hd__buf_2 fanout204 (.A(net827),
    .X(net826));
 sky130_fd_sc_hd__buf_8 fanout205 (.A(net828),
    .X(net827));
 sky130_fd_sc_hd__buf_6 fanout206 (.A(net730),
    .X(net828));
 sky130_fd_sc_hd__clkbuf_4 fanout207 (.A(net830),
    .X(net829));
 sky130_fd_sc_hd__buf_2 fanout208 (.A(net31),
    .X(net830));
 sky130_fd_sc_hd__buf_2 fanout209 (.A(net833),
    .X(net831));
 sky130_fd_sc_hd__clkbuf_4 fanout210 (.A(net833),
    .X(net832));
 sky130_fd_sc_hd__buf_2 fanout211 (.A(net834),
    .X(net833));
 sky130_fd_sc_hd__buf_2 fanout212 (.A(net31),
    .X(net834));
 sky130_fd_sc_hd__buf_4 wire213 (.A(net22),
    .X(net835));
 sky130_fd_sc_hd__buf_8 max_cap214 (.A(net17),
    .X(net836));
 sky130_fd_sc_hd__buf_4 fanout215 (.A(net838),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_8 fanout216 (.A(net839),
    .X(net838));
 sky130_fd_sc_hd__buf_8 fanout217 (.A(net16),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_4 fanout218 (.A(net791),
    .X(net840));
 sky130_fd_sc_hd__clkbuf_8 fanout219 (.A(net801),
    .X(net841));
 sky130_fd_sc_hd__buf_4 fanout220 (.A(net602),
    .X(net842));
 sky130_fd_sc_hd__buf_4 fanout221 (.A(net753),
    .X(net843));
 sky130_fd_sc_hd__clkbuf_4 fanout222 (.A(net601),
    .X(net844));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout223 (.A(net601),
    .X(net845));
 sky130_fd_sc_hd__buf_4 fanout224 (.A(net572),
    .X(net846));
 sky130_fd_sc_hd__buf_4 fanout225 (.A(net701),
    .X(net847));
 sky130_fd_sc_hd__buf_4 fanout226 (.A(net849),
    .X(net848));
 sky130_fd_sc_hd__buf_4 fanout227 (.A(net627),
    .X(net849));
 sky130_fd_sc_hd__buf_4 fanout228 (.A(net665),
    .X(net850));
 sky130_fd_sc_hd__clkbuf_8 fanout229 (.A(net624),
    .X(net851));
 sky130_fd_sc_hd__buf_12 fanout230 (.A(net182),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net615 (.A(net615),
    .X(clknet_0_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net615 (.A(clknet_0_net615),
    .X(clknet_1_0__leaf_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net615 (.A(clknet_0_net615),
    .X(clknet_1_1__leaf_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net475 (.A(net475),
    .X(clknet_0_net475));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net475 (.A(clknet_0_net475),
    .X(clknet_1_0__leaf_net475));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net475 (.A(clknet_0_net475),
    .X(clknet_1_1__leaf_net475));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net799 (.A(net799),
    .X(clknet_0_net799));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net799 (.A(clknet_0_net799),
    .X(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net799 (.A(clknet_0_net799),
    .X(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net370 (.A(net370),
    .X(clknet_0_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net370 (.A(clknet_0_net370),
    .X(clknet_1_0__leaf_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net370 (.A(clknet_0_net370),
    .X(clknet_1_1__leaf_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net512 (.A(net512),
    .X(clknet_0_net512));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net512 (.A(clknet_0_net512),
    .X(clknet_1_0__leaf_net512));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net512 (.A(clknet_0_net512),
    .X(clknet_1_1__leaf_net512));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net295 (.A(net295),
    .X(clknet_0_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net295 (.A(clknet_0_net295),
    .X(clknet_1_0__leaf_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net295 (.A(clknet_0_net295),
    .X(clknet_1_1__leaf_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net400 (.A(net400),
    .X(clknet_0_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net400 (.A(clknet_0_net400),
    .X(clknet_1_0__leaf_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net400 (.A(clknet_0_net400),
    .X(clknet_1_1__leaf_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net300 (.A(net300),
    .X(clknet_0_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net300 (.A(clknet_0_net300),
    .X(clknet_1_0__leaf_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net300 (.A(clknet_0_net300),
    .X(clknet_1_1__leaf_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net289 (.A(net289),
    .X(clknet_0_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net289 (.A(clknet_0_net289),
    .X(clknet_1_0__leaf_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net289 (.A(clknet_0_net289),
    .X(clknet_1_1__leaf_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net305 (.A(net305),
    .X(clknet_0_net305));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net305 (.A(clknet_0_net305),
    .X(clknet_1_0__leaf_net305));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net305 (.A(clknet_0_net305),
    .X(clknet_1_1__leaf_net305));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net301 (.A(net301),
    .X(clknet_0_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net301 (.A(clknet_0_net301),
    .X(clknet_1_0__leaf_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net301 (.A(clknet_0_net301),
    .X(clknet_1_1__leaf_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net268 (.A(net268),
    .X(clknet_0_net268));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net268 (.A(clknet_0_net268),
    .X(clknet_1_0__leaf_net268));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net268 (.A(clknet_0_net268),
    .X(clknet_1_1__leaf_net268));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net255 (.A(net255),
    .X(clknet_0_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net255 (.A(clknet_0_net255),
    .X(clknet_1_0__leaf_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net255 (.A(clknet_0_net255),
    .X(clknet_1_1__leaf_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net614 (.A(net614),
    .X(clknet_0_net614));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net614 (.A(clknet_0_net614),
    .X(clknet_1_0__leaf_net614));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net614 (.A(clknet_0_net614),
    .X(clknet_1_1__leaf_net614));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net473 (.A(net473),
    .X(clknet_0_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net473 (.A(clknet_0_net473),
    .X(clknet_1_0__leaf_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net473 (.A(clknet_0_net473),
    .X(clknet_1_1__leaf_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net793 (.A(net793),
    .X(clknet_0_net793));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net793 (.A(clknet_0_net793),
    .X(clknet_1_0__leaf_net793));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net793 (.A(clknet_0_net793),
    .X(clknet_1_1__leaf_net793));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net367 (.A(net367),
    .X(clknet_0_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net367 (.A(clknet_0_net367),
    .X(clknet_1_0__leaf_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net367 (.A(clknet_0_net367),
    .X(clknet_1_1__leaf_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net198 (.A(net198),
    .X(clknet_0_net198));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net198 (.A(clknet_0_net198),
    .X(clknet_1_0__leaf_net198));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net198 (.A(clknet_0_net198),
    .X(clknet_1_1__leaf_net198));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net199 (.A(net199),
    .X(clknet_0_net199));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net199 (.A(clknet_0_net199),
    .X(clknet_1_0__leaf_net199));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net199 (.A(clknet_0_net199),
    .X(clknet_1_1__leaf_net199));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net200 (.A(net200),
    .X(clknet_0_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net200 (.A(clknet_0_net200),
    .X(clknet_1_0__leaf_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net200 (.A(clknet_0_net200),
    .X(clknet_1_1__leaf_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net179 (.A(net179),
    .X(clknet_0_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_0__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_1__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net178 (.A(net178),
    .X(clknet_0_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net178 (.A(clknet_0_net178),
    .X(clknet_1_0__leaf_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net178 (.A(clknet_0_net178),
    .X(clknet_1_1__leaf_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net375 (.A(net375),
    .X(clknet_0_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net375 (.A(clknet_0_net375),
    .X(clknet_1_0__leaf_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net375 (.A(clknet_0_net375),
    .X(clknet_1_1__leaf_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net277 (.A(net277),
    .X(clknet_0_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net277 (.A(clknet_0_net277),
    .X(clknet_1_0__leaf_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net277 (.A(clknet_0_net277),
    .X(clknet_1_1__leaf_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net281 (.A(net281),
    .X(clknet_0_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net281 (.A(clknet_0_net281),
    .X(clknet_1_0__leaf_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net281 (.A(clknet_0_net281),
    .X(clknet_1_1__leaf_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net282 (.A(net282),
    .X(clknet_0_net282));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net282 (.A(clknet_0_net282),
    .X(clknet_1_0__leaf_net282));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net282 (.A(clknet_0_net282),
    .X(clknet_1_1__leaf_net282));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net276 (.A(net276),
    .X(clknet_0_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net276 (.A(clknet_0_net276),
    .X(clknet_1_0__leaf_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net276 (.A(clknet_0_net276),
    .X(clknet_1_1__leaf_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net166 (.A(net166),
    .X(clknet_0_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net166 (.A(clknet_0_net166),
    .X(clknet_1_0__leaf_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net166 (.A(clknet_0_net166),
    .X(clknet_1_1__leaf_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net769 (.A(net769),
    .X(clknet_0_net769));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net769 (.A(clknet_0_net769),
    .X(clknet_1_0__leaf_net769));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net769 (.A(clknet_0_net769),
    .X(clknet_1_1__leaf_net769));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net162 (.A(net162),
    .X(clknet_0_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net162 (.A(clknet_0_net162),
    .X(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net162 (.A(clknet_0_net162),
    .X(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net161 (.A(net161),
    .X(clknet_0_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net161 (.A(clknet_0_net161),
    .X(clknet_1_0__leaf_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net161 (.A(clknet_0_net161),
    .X(clknet_1_1__leaf_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net159 (.A(net159),
    .X(clknet_0_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net159 (.A(clknet_0_net159),
    .X(clknet_1_0__leaf_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net159 (.A(clknet_0_net159),
    .X(clknet_1_1__leaf_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net766 (.A(net766),
    .X(clknet_0_net766));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net766 (.A(clknet_0_net766),
    .X(clknet_1_0__leaf_net766));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net766 (.A(clknet_0_net766),
    .X(clknet_1_1__leaf_net766));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net786 (.A(net786),
    .X(clknet_0_net786));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net786 (.A(clknet_0_net786),
    .X(clknet_1_0__leaf_net786));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net786 (.A(clknet_0_net786),
    .X(clknet_1_1__leaf_net786));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net742 (.A(net742),
    .X(clknet_0_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net742 (.A(clknet_0_net742),
    .X(clknet_1_0__leaf_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net742 (.A(clknet_0_net742),
    .X(clknet_1_1__leaf_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net97 (.A(net97),
    .X(clknet_0_net97));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net97 (.A(clknet_0_net97),
    .X(clknet_1_0__leaf_net97));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net97 (.A(clknet_0_net97),
    .X(clknet_1_1__leaf_net97));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net800 (.A(net800),
    .X(clknet_0_net800));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net800 (.A(clknet_0_net800),
    .X(clknet_1_0__leaf_net800));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net800 (.A(clknet_0_net800),
    .X(clknet_1_1__leaf_net800));
 sky130_fd_sc_hd__buf_2 rebuffer1 (.A(net771),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net903),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net903),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_1 rebuffer4 (.A(net855),
    .X(net856));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer5 (.A(net856),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net46),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net858),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net125),
    .X(net860));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer9 (.A(net860),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net861),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net861),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net57),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net57),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net732),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net803),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net828),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net868),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net828),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net870),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net871),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net872),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net740),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net728),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net875),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net876),
    .X(net877));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer26 (.A(net139),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(net878),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(net878),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net228),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(net228),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer31 (.A(net882),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(net813),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(net884),
    .X(net885));
 sky130_fd_sc_hd__clkbuf_4 clone34 (.A(net740),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer35 (.A(net21),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer36 (.A(net887),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer37 (.A(net890),
    .X(net889));
 sky130_fd_sc_hd__clkbuf_1 clone38 (.A(net182),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer39 (.A(net43),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer40 (.A(net891),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net608),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net429),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net572),
    .X(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in62));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in63));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in64));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(in65));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(in66));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(in67));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(in68));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(in69));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(in70));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(in71));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(in72));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(in73));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(in74));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(in75));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(in76));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(in77));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(in78));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(in79));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(in80));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(in81));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(in82));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(in83));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(in84));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(in85));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(in86));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(in87));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(in88));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(in89));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(in90));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(in91));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(in92));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(in93));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(in94));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(in95));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(in96));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(in97));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(in98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(in99));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_X (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_Y (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S0 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_Y (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A3 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A3 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_X (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A3 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_X (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A0 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A3 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A3 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A3 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_Y (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A0 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_Y (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A4 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_D (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_S1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A0 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_B1_N (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_X (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_Y (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A4 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A3 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_Y (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A4 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A3 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A3 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_X (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A0 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A3 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A0 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A3 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_X (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A3 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A3 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_X (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_SCD (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_X (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_S1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_X (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A4 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_B1_N (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_X (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_B1_N (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_Y (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A3 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A4 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A3 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_B1_N (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_X (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer26_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A2 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_B1_N (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_X (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_X (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S0 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A3 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A4 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_X (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A0 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A4 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A3 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_X (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A0 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A0 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_X (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A3 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A0 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A0 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_X (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A0 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_X (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A3 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_X (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_S0 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A0 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_S0 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S0 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S0 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A4 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_X (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_X (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A3 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_X (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_A3 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_X (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A0 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A3 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_X (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_B1_N (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_Y (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_S1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A0 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A0 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_X (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A3 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S0 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A3 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_X (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_X (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_S0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_X (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_B1_N (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_X (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_X (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S0 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A4 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_X (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_X (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S0 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_B1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_X (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_X (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A0 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_B1_N (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_Y (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A3 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_Y (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B1_N (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_B1_N (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_B1_N (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A3 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_X (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_S0 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_A3 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_X (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A3 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A4 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_B1_N (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_Y (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_B1_N (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_X (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire213_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A3 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_Y (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A3 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A0 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_B1_N (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A2 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S0 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A2 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_X (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A4 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_X (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A3 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_X (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A0 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A0 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A4 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A3 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_X (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A3 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A3 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A0 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_B1_N (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_X (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A2 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S0 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A3 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A3 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_B1_N (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_X (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A3 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A2 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_S0 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_X (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_S0 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_X (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A3 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_B1_N (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_S0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_X (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_S0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_X (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A0 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A4 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_X (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A2 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_X (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_X (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A4 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S0 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_X (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A3 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A2 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_B1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S0 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A2 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_X (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A3 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_X (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S0 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_X (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_X (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_B1_N (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A2 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A2 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_B1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A3 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S0 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_X (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A3 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_X (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A3 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_X (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_X (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A0 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A3 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_B (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_X (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_B1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_Y (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A3 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S0 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_X (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A0 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A4 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A4 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_B1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_X (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S0 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A3 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_B1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_Y (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A3 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_S0 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_X (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A0 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_S0 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_B1_N (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A3 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A4 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A3 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_X (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_Y (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A0 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_X (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_B1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_B1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_B1_N (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_B1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A4 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_X (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A0 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A2 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_B1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A3 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_X (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_X (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A4 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A3 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A2 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_X (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_D (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A3 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_X (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A0 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A3 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A3 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A2 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A3 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A2 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_SCE (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_X (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A2 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A2 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_Q (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A3 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A0 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A3 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A4 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_X (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_B1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_X (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A0 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A3 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A3 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_X (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A3 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_X (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_D (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_X (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_X (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_X (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A3 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A1 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A3 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_X (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_X (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_X (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_X (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_B (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_X (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_B1_N (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_X (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A2 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A2 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A2 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_X (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A0 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A2 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S0 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_X (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A0 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A3 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A3 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A3 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_SCE (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_X (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A3 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_X (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A2 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A4 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_SCD (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_SCE (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A3 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_X (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold42_A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A3 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_Q (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer39_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A3 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_S0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A3 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A3 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_X (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A0 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A2 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_X (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A2 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A3 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A3 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_X (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_D (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_X (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A4 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_X (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A0 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_X (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A2 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S0 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A2 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_X (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A0 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A3 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A3 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_B1_N (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_B1_N (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_X (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_B1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_X (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_X (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_X (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A3 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_S1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_X (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A0 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A4 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_B1_N (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_X (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A3 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_B1_N (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_S0 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S0 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_X (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_Q (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S0 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_B1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A0 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B1_N (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_X (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_D (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_Y (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge877_D (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_Y (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A3 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_B1_N (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A0 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A4 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_X (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_Q (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_S0 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S0 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S0 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S0 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_Q (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A3 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S0 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_B1 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_B1 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_Q_N (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_Q (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A4 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_B1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_B1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_S1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_Q_N (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S1 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold41_A (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_Q (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S0 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S0 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_S1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_B1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_Q (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_S1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_S1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A3 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_X (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge877_Q (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S0 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_S0 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S0 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_B1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_S0 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_Q_N (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_Q (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S1 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S1 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S1 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S1 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_B1 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_Q_N (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_S1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A3 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_S1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_Q (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_S1 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_S1 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S0 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_Q (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_S0 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A3 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A3 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_X (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S0 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_B1_N (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A3 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A3 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_X (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_B1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A3 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_B1_N (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_X (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_X (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A3 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B1_N (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A3 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_X (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A3 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_X (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A3 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A3 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A3 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A3 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_X (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_X (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_S0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_S1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_S1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A3 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_X (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_X (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone38_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A3 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_A (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A1 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A3 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A3 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A0 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S0 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A4 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A3 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_B1_N (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A4 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A0 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A4 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_B (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A3 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A0 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A0 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B1_N (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A0 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A2 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A0 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A3 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A1 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A2 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A0 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B1_N (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A2 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A1 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A3 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A0 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A2 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A1 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A3 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A2 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A2 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A1 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_S0 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A1 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A1 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A2 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A1 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A2 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A1 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A2 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A2 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A2 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_B1_N (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_B (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A2 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A0 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A4 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A3 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A1 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A3 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_B1 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_S0 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B1_N (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A1 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A0 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A3 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A3 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A2 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A2 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A4 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A3 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_B1_N (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A2 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A2 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_B1_N (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A3 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A1 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B1 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A2 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B1_N (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A3 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A1 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A2 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A1 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A2 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A2 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A3 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A0 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A2 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S0 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A2 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A0 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S0 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A1 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S0 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A4 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_X (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A0 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A2 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A2 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_B1 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A1 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S0 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A3 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_B1_N (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B1_N (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A1 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A1 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A3 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_S0 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B1_N (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A1 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_B1_N (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A1 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A3 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A0 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_B1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S1 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A3 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A2 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A1 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A3 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A0 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_S0 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A3 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S0 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A2 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_SET_B (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A1 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A1 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A2 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A2 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A2 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A3 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_RESET_B (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_B1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_S1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_X (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A2 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S1 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A3 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A2 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A2 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_S1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_B1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_A (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A2 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_S1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A2 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_X (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A2 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A3 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_S0 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_B1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A3 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A0 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A2 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A3 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A3 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A3 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A3 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A0 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A0 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_B1_N (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_B1_N (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A4 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A0 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_B1_N (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A2 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A2 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A3 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A0 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A2 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A2 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A2 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_X (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A2 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A3 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A2 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A3 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A1 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A0 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A4 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_B1_N (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A0 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S0 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A4 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_X (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A0 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A1 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A1 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S1 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A0 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A0 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A3 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A2 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_S1 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A1 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A3 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A3 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A2 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A1 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_B1_N (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A2 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_A2 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_X (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A0 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S0 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A4 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A2 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A1 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A2 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A3 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_X (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A3 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A3 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_B1_N (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_X (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A3 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A0 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A0 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A4 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_B1_N (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A3 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_X (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_X (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_X (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A3 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A2 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A2 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_S0 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_B1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A2 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_X (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A3 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A0 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A2 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A2 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A3 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_X (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A0 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A2 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A4 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_X (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S0 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A1 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_S1 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_B1_N (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_X (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A2 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A1 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A3 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_B1_N (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_X (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A1 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A3 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A2 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A2 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_X (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_S1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A2 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A2 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_X (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A2 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A3 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A3 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_A1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_X (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A0 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A3 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_X (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A1 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A1 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_X (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A0 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S0 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A2 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A2 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_X (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_B1_N (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A2 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_S0 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_B (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_X (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A0 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A2 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_X (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A3 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A4 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_X (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A3 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S0 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A2 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_X (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A3 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A3 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A4 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_X (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A1 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A3 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A3 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_X (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A1 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A1 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A2 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A2 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A2 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A3 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A1 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A2 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A4 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_B1 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_X (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A2 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A4 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A4 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_X (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A3 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A1 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_S1 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_X (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A2 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_B1_N (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_X (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A2 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A1 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A2 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_X (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A0 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A4 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A4 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A2 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_X (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A3 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S0 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A3 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_B1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_B1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S0 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A3 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S0 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A3 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A2 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A2 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A2 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_B1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_X (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_S0 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A3 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A3 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A2 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_X (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S0 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A3 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_X (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A4 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_B (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A3 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_Y (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_X (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A2 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A2 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A3 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A3 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_X (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer14_A (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_X (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_Q_N (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S0 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S0 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S0 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_B1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A4 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_X (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A1 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_X (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S0 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A2 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_X (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A3 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A2 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A3 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S0 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_X (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_X (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone34_A (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer22_A (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_Q (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S0 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S0 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_S1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_B1_N (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_B1_N (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap201_A (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S1 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S0 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A3 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_B1 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_X (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A2 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A2 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A0 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_X (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_S0 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_SCD (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_X (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S0 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_X (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A3 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_X (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_output129_A (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_X (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_output130_A (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S0 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A3 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A2 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_X (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_Q (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_B1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A1 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A3 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A0 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_X (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_output133_A (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_S0 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A2 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_X (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_output134_A (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A4 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_B1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_X (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_S0 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S0 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A4 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A2 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A3 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_B1_N (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_B1_N (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_X (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_output136_A (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A2 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A4 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_X (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_output137_A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_Q (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S0 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_S0 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A2 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A2 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A3 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A0 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A2 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_X (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_output139_A (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A2 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_S1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A2 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B1_N (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_X (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_output140_A (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S0 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A2 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_X (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_output141_A (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A3 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_X (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_A (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A1 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A1 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_X (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_output145_A (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_S1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A2 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_B1_N (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_B1_N (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_X (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_output148_A (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A3 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A4 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A3 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_X (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer3_A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A3 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_output151_A (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A2 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_X (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_output155_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_S0 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A2 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B1_N (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A0 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_output157_A (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A1 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A3 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_X (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_output158_A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A3 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A2 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_X (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_output161_A (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S0 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A2 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_S0 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_X (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_output163_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_X (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_output165_A (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A2 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_X (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_S0 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_S1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_Y (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_output174_A (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A3 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_X (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_output175_A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A2 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A3 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A4 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_X (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_A (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_output179_A (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_Q (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S0 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S0 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S0 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_X (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_B1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A3 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S0 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A3 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B1_N (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_X (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_X (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A3 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_B1_N (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_X (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_S0 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A3 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A4 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A0 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A3 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_S0 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A2 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A4 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_B1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_X (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_B1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A3 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A3 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A2 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A3 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A4 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_X (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A3 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A2 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A3 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A2 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A2 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_B1_N (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A4 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_S1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_B (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_X (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A4 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A2 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_B1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A4 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_S0 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A2 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A3 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A3 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_X (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A2 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S0 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_B1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A2 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A4 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A4 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_B1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_B1_N (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_X (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A2 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer32_A (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_X (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A2 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A2 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A3 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_B1_N (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_B1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_X (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_B1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A3 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A3 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B1_N (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_B1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_B1_N (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A4 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A3 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap193_X (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A2 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S0 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_X (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A3 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S0 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A2 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A3 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A3 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_X (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A4 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A3 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_B1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_X (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S0 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A1 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A2 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_B1_N (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A4 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_X (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A3 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A3 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_B1_N (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A3 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B1_N (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap198_X (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A3 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_X (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_S1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_B1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_B1_N (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_B1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_B1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_B1_N (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A2 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_X (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_B1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap201_X (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_SET_B (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_X (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A3 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_S1 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_B1_N (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_B1_N (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A1 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_S0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_RESET_B (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A2 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_B1 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_X (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_S0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_S0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B1_N (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_B1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_B1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_B1_N (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_B1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_B1_N (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_B1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_X (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B1_N (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_B1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_B1_N (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_S1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_X (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_S0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_B1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer18_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer16_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_X (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A3 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_B1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_X (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B1_N (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A3 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_B1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_S1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_B1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_SET_B (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_B1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_B1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_S1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A2 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_X (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_B1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A3 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_X (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B1_N (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_B1_N (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A3 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A3 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A2 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B1_N (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_B1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_S1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_X (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_B1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_B1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_S1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_B1_N (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A4 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_B1_N (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A4 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_X (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A3 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A4 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_B1_N (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_B1_N (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_X (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_B1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_B1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_B1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire213_X (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A2 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A3 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_X (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B1_N (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A4 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_S0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_B1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_B1_N (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_B1_N (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_X (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_B1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A3 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_B1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A4 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_B1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A4 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A3 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_S0 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_X (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A3 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_B1_N (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_A3 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_B1_N (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_B1_N (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_B (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_B (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_output169_A (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_X (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_S1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_B1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_X (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_B1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A3 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_B1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_B1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_X (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_B1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_B1_N (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_A (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A3 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_S0 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_X (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_B1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_B1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A4 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_X (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A4 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_B1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_B1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_B1_N (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_B1_N (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S0 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_S0 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_S1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_B1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A2 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_X (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S0 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_S0 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_SCE (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_B1_N (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A3 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B1_N (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_X (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_B1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_B1_N (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S0 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A2 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_X (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A2 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_B1_N (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_B1_N (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B1_N (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_X (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_S0 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A3 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A3 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A0 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S0 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A3 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A3 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S1 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A2 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_X (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A2 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S0 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S0 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S0 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_S0 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A3 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A2 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_X (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A2 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B1_N (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_CLK_N (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_CLK_N (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_CLK_N (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_CLK_N (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_CLK_N (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_GATE (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_X (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_GATE (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_GATE_N (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge877_GATE (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_X (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_GATE_N (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_GATE_N (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_GATE (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge875_GATE (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_X (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_GATE_N (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_GATE_N (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_X (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_B1 (.DIODE(clknet_1_0__leaf_net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S1 (.DIODE(clknet_1_0__leaf_net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S1 (.DIODE(clknet_1_0__leaf_net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A3 (.DIODE(clknet_1_0__leaf_net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net615_X (.DIODE(clknet_1_0__leaf_net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_S1 (.DIODE(clknet_1_1__leaf_net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S0 (.DIODE(clknet_1_1__leaf_net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S1 (.DIODE(clknet_1_1__leaf_net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_S0 (.DIODE(clknet_1_1__leaf_net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net615_X (.DIODE(clknet_1_1__leaf_net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_B1 (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S1 (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_B1 (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_B1 (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S1 (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_S1 (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S1 (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S1 (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net799_X (.DIODE(clknet_1_0__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_S1 (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_B1 (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_B1_N (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S1 (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_B1 (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_B1_N (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S1 (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_B1 (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_B1_N (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S1 (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_output177_A (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net799_X (.DIODE(clknet_1_1__leaf_net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_B1_N (.DIODE(clknet_1_0__leaf_net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S1 (.DIODE(clknet_1_0__leaf_net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_S1 (.DIODE(clknet_1_0__leaf_net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_B1 (.DIODE(clknet_1_0__leaf_net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_B1 (.DIODE(clknet_1_0__leaf_net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net614_X (.DIODE(clknet_1_0__leaf_net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_S1 (.DIODE(clknet_1_1__leaf_net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S1 (.DIODE(clknet_1_1__leaf_net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net614_X (.DIODE(clknet_1_1__leaf_net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A1 (.DIODE(clknet_1_0__leaf_net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A4 (.DIODE(clknet_1_0__leaf_net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net769_X (.DIODE(clknet_1_0__leaf_net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net162_A (.DIODE(clknet_0_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net162_A (.DIODE(clknet_0_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net162_X (.DIODE(clknet_0_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A3 (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_B1 (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S0 (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_SCD (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A1 (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A0 (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net162_X (.DIODE(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S0 (.DIODE(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A3 (.DIODE(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_B1 (.DIODE(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A3 (.DIODE(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A1 (.DIODE(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_A0 (.DIODE(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net162_X (.DIODE(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_B1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer6_X (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer17_A (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer16_X (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer22_X (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer25_A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_S0 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer24_X (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer28_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer27_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A4 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer26_X (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A3 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer33_A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer32_X (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer33_X (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone34_X (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_S1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer37_X (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_B1_N (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A4 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer37_A (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone38_X (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net653));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(net53),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer38 (.A(net896),
    .X(net897));
 sky130_fd_sc_hd__mux4_1 clone39 (.A0(net21),
    .A1(net28),
    .A2(net818),
    .A3(net823),
    .S0(net904),
    .S1(net903),
    .X(net898));
 sky130_fd_sc_hd__mux4_1 clone40 (.A0(net20),
    .A1(net820),
    .A2(net712),
    .A3(net633),
    .S0(net825),
    .S1(net837),
    .X(net899));
 sky130_fd_sc_hd__a21bo_1 clone41 (.A1(net847),
    .A2(net21),
    .B1_N(net838),
    .X(net900));
 sky130_fd_sc_hd__a21bo_1 clone42 (.A1(net760),
    .A2(net630),
    .B1_N(net849),
    .X(net901));
 sky130_fd_sc_hd__mux4_1 clone43 (.A0(net21),
    .A1(net28),
    .A2(net818),
    .A3(net823),
    .S0(net904),
    .S1(net771),
    .X(net902));
 sky130_fd_sc_hd__mux4_1 clone44 (.A0(net20),
    .A1(net820),
    .A2(net712),
    .A3(net633),
    .S0(net825),
    .S1(net837),
    .X(net903));
 sky130_fd_sc_hd__a21bo_1 clone45 (.A1(net760),
    .A2(net630),
    .B1_N(net849),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer46 (.A(net463),
    .X(net905));
 sky130_fd_sc_hd__a21bo_1 clone47 (.A1(net837),
    .A2(net18),
    .B1_N(net632),
    .X(net906));
 sky130_fd_sc_hd__a21bo_1 clone48 (.A1(net131),
    .A2(net908),
    .B1_N(net642),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer49 (.A(net136),
    .X(net908));
 sky130_fd_sc_hd__clkbuf_1 clone50 (.A(net740),
    .X(net909));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
