module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in3,
    in4,
    in5,
    in6,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out3,
    out4,
    out5,
    out6,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in3;
 input in4;
 input in5;
 input in6;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out3;
 output out4;
 output out5;
 output out6;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_0_net390;
 wire clknet_1_0__leaf_net390;
 wire clknet_1_1__leaf_net390;
 wire clknet_0_net757;
 wire clknet_1_0__leaf_net757;
 wire clknet_1_1__leaf_net757;
 wire clknet_0_net814;
 wire clknet_1_0__leaf_net814;
 wire clknet_1_1__leaf_net814;
 wire clknet_0_net596;
 wire clknet_1_0__leaf_net596;
 wire clknet_1_1__leaf_net596;
 wire clknet_0_net432;
 wire clknet_1_0__leaf_net432;
 wire clknet_1_1__leaf_net432;
 wire clknet_0_net463;
 wire clknet_1_0__leaf_net463;
 wire clknet_1_1__leaf_net463;
 wire clknet_0_net261;
 wire clknet_1_0__leaf_net261;
 wire clknet_1_1__leaf_net261;
 wire clknet_0_net399;
 wire clknet_1_0__leaf_net399;
 wire clknet_1_1__leaf_net399;
 wire clknet_0_net402;
 wire clknet_1_0__leaf_net402;
 wire clknet_1_1__leaf_net402;
 wire clknet_0_net398;
 wire clknet_1_0__leaf_net398;
 wire clknet_1_1__leaf_net398;
 wire clknet_0_net401;
 wire clknet_1_0__leaf_net401;
 wire clknet_1_1__leaf_net401;
 wire clknet_0_net250;
 wire clknet_1_0__leaf_net250;
 wire clknet_1_1__leaf_net250;
 wire clknet_0_net287;
 wire clknet_1_0__leaf_net287;
 wire clknet_1_1__leaf_net287;
 wire clknet_0_net449;
 wire clknet_1_0__leaf_net449;
 wire clknet_1_1__leaf_net449;
 wire clknet_0_net258;
 wire clknet_1_0__leaf_net258;
 wire clknet_1_1__leaf_net258;
 wire clknet_0_net252;
 wire clknet_1_0__leaf_net252;
 wire clknet_1_1__leaf_net252;
 wire clknet_0_net539;
 wire clknet_1_0__leaf_net539;
 wire clknet_1_1__leaf_net539;
 wire clknet_0_net253;
 wire clknet_1_0__leaf_net253;
 wire clknet_1_1__leaf_net253;
 wire clknet_0_net517;
 wire clknet_1_0__leaf_net517;
 wire clknet_1_1__leaf_net517;
 wire clknet_0_net255;
 wire clknet_1_0__leaf_net255;
 wire clknet_1_1__leaf_net255;
 wire clknet_0_net251;
 wire clknet_1_0__leaf_net251;
 wire clknet_1_1__leaf_net251;
 wire clknet_0_net290;
 wire clknet_1_0__leaf_net290;
 wire clknet_1_1__leaf_net290;
 wire clknet_0_net260;
 wire clknet_1_0__leaf_net260;
 wire clknet_1_1__leaf_net260;
 wire clknet_0_net242;
 wire clknet_1_0__leaf_net242;
 wire clknet_1_1__leaf_net242;
 wire clknet_0_net356;
 wire clknet_1_0__leaf_net356;
 wire clknet_1_1__leaf_net356;
 wire clknet_0_net359;
 wire clknet_1_0__leaf_net359;
 wire clknet_1_1__leaf_net359;
 wire clknet_0_net160;
 wire clknet_1_0__leaf_net160;
 wire clknet_1_1__leaf_net160;
 wire clknet_0_net165;
 wire clknet_1_0__leaf_net165;
 wire clknet_1_1__leaf_net165;
 wire clknet_0_net294;
 wire clknet_1_0__leaf_net294;
 wire clknet_1_1__leaf_net294;
 wire clknet_0_net166;
 wire clknet_1_0__leaf_net166;
 wire clknet_1_1__leaf_net166;
 wire clknet_0_net158;
 wire clknet_1_0__leaf_net158;
 wire clknet_1_1__leaf_net158;
 wire clknet_0_net171;
 wire clknet_1_0__leaf_net171;
 wire clknet_1_1__leaf_net171;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;

 sky130_fd_sc_hd__and2_2 c100 (.A(net79),
    .B(net44),
    .X(net82));
 sky130_fd_sc_hd__sdfxtp_2 c101 (.CLK(clknet_leaf_28_clk),
    .D(net68),
    .SCD(net81),
    .SCE(net79),
    .Q(net83));
 sky130_fd_sc_hd__mux4_1 c102 (.A0(net66),
    .A1(net80),
    .A2(net77),
    .A3(net82),
    .S0(net83),
    .S1(net63),
    .X(net84));
 sky130_fd_sc_hd__and2_1 c103 (.A(net81),
    .B(net83),
    .X(net85));
 sky130_fd_sc_hd__sdfxtp_1 c104 (.CLK(clknet_leaf_27_clk),
    .D(net80),
    .SCD(net36),
    .SCE(net856),
    .Q(net86));
 sky130_fd_sc_hd__clkbuf_1 c105 (.A(net4),
    .X(net87));
 sky130_fd_sc_hd__sdfxtp_1 c106 (.CLK(clknet_leaf_28_clk),
    .D(net949),
    .SCD(net10),
    .SCE(net80),
    .Q(net88));
 sky130_fd_sc_hd__clkbuf_1 c107 (.A(net48),
    .X(net89));
 sky130_fd_sc_hd__and2_0 c108 (.A(net71),
    .B(net942),
    .X(net90));
 sky130_fd_sc_hd__dfbbn_1 c109 (.CLK_N(clknet_leaf_28_clk),
    .D(net90),
    .RESET_B(net68),
    .SET_B(net74),
    .Q(net91));
 sky130_fd_sc_hd__clkbuf_1 c110 (.A(net736),
    .X(net92));
 sky130_fd_sc_hd__buf_1 c111 (.A(net91),
    .X(net93));
 sky130_fd_sc_hd__buf_1 c112 (.A(net65),
    .X(net94));
 sky130_fd_sc_hd__buf_1 c113 (.A(net89),
    .X(net95));
 sky130_fd_sc_hd__and2_0 c114 (.A(net92),
    .B(net804),
    .X(net96));
 sky130_fd_sc_hd__and3_1 c115 (.A(net94),
    .B(net85),
    .C(net21),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_1 c116 (.A(net735),
    .X(net97));
 sky130_fd_sc_hd__or4bb_2 c117 (.A(net95),
    .B(net97),
    .C_N(net93),
    .D_N(net8),
    .X(net98));
 sky130_fd_sc_hd__and2_1 c118 (.A(net21),
    .B(net88),
    .X(net99));
 sky130_fd_sc_hd__dlrbn_1 c119 (.D(net98),
    .GATE_N(clknet_leaf_26_clk),
    .RESET_B(net93),
    .Q(net100));
 sky130_fd_sc_hd__dlrbn_1 c120 (.D(net87),
    .GATE_N(clknet_leaf_26_clk),
    .RESET_B(net94),
    .Q(net824),
    .Q_N(net101));
 sky130_fd_sc_hd__buf_1 c121 (.A(net96),
    .X(net826));
 sky130_fd_sc_hd__dlrbp_1 c122 (.D(net868),
    .GATE(clknet_leaf_26_clk),
    .RESET_B(net98),
    .Q(net810),
    .Q_N(net102));
 sky130_fd_sc_hd__dfbbn_1 c123 (.CLK_N(clknet_leaf_28_clk),
    .D(net97),
    .RESET_B(net826),
    .SET_B(net87),
    .Q(net103));
 sky130_fd_sc_hd__and2_0 c124 (.A(net103),
    .B(net101),
    .X(net104));
 sky130_fd_sc_hd__and2_0 c125 (.A(net10),
    .B(net826),
    .X(net105));
 sky130_fd_sc_hd__dlymetal6s2s_1 c126 (.A(net806),
    .X(net106));
 sky130_fd_sc_hd__and2_2 c127 (.A(net804),
    .B(net106),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 c128 (.A(net786),
    .X(net108));
 sky130_fd_sc_hd__and2_1 c129 (.A(net792),
    .B(net808),
    .X(net109));
 sky130_fd_sc_hd__and2_2 c130 (.A(net805),
    .B(net786),
    .X(net110));
 sky130_fd_sc_hd__and2_2 c131 (.A(net108),
    .B(net107),
    .X(net111));
 sky130_fd_sc_hd__and2_2 c132 (.A(net793),
    .B(net107),
    .X(net112));
 sky130_fd_sc_hd__buf_1 c133 (.A(net733),
    .X(net113));
 sky130_fd_sc_hd__buf_1 c134 (.A(net107),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 c135 (.A(net733),
    .X(net115));
 sky130_fd_sc_hd__dlrbp_1 c136 (.D(net113),
    .GATE(clknet_leaf_2_clk),
    .RESET_B(net111),
    .Q(net117),
    .Q_N(net116));
 sky130_fd_sc_hd__dlrtn_1 c137 (.D(net794),
    .GATE_N(clknet_leaf_3_clk),
    .RESET_B(net114),
    .Q(net118));
 sky130_fd_sc_hd__dlrtn_1 c138 (.D(net106),
    .GATE_N(clknet_leaf_2_clk),
    .RESET_B(net112),
    .Q(net119));
 sky130_fd_sc_hd__dlrtn_1 c139 (.D(net114),
    .GATE_N(clknet_leaf_3_clk),
    .RESET_B(net109),
    .Q(net120));
 sky130_fd_sc_hd__and2_4 c140 (.A(net109),
    .B(net107),
    .X(net121));
 sky130_fd_sc_hd__dlrtp_1 c141 (.D(net111),
    .GATE(clknet_leaf_2_clk),
    .RESET_B(net914),
    .Q(net122));
 sky130_fd_sc_hd__and2_1 c142 (.A(net120),
    .B(net794),
    .X(net123));
 sky130_fd_sc_hd__and2_1 c143 (.A(net115),
    .B(net123),
    .X(net124));
 sky130_fd_sc_hd__mux4_1 c144 (.A0(net792),
    .A1(net118),
    .A2(net122),
    .A3(net121),
    .S0(net111),
    .S1(net115),
    .X(net125));
 sky130_fd_sc_hd__and2_2 c145 (.A(net124),
    .B(net123),
    .X(net126));
 sky130_fd_sc_hd__and2_1 c146 (.A(net802),
    .B(net124),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 c147 (.A(net753),
    .X(net128));
 sky130_fd_sc_hd__buf_1 c148 (.A(in10),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 c149 (.A(net752),
    .X(net130));
 sky130_fd_sc_hd__and2_1 c150 (.A(net4),
    .B(net113),
    .X(net131));
 sky130_fd_sc_hd__dlrtp_1 c151 (.D(net7),
    .GATE(clknet_leaf_38_clk),
    .RESET_B(net131),
    .Q(net132));
 sky130_fd_sc_hd__and2_1 c152 (.A(net7),
    .B(net756),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 c153 (.A(net956),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_4 c154 (.A(net128),
    .X(net830));
 sky130_fd_sc_hd__and2_2 c155 (.A(net133),
    .B(net129),
    .X(net135));
 sky130_fd_sc_hd__dlrtp_1 c156 (.D(net16),
    .GATE(clknet_leaf_38_clk),
    .RESET_B(net111),
    .Q(net136));
 sky130_fd_sc_hd__and2_0 c157 (.A(net118),
    .B(net110),
    .X(net137));
 sky130_fd_sc_hd__and3_4 c158 (.A(net802),
    .B(net7),
    .C(net119),
    .X(net138));
 sky130_fd_sc_hd__and3_1 c159 (.A(net134),
    .B(net960),
    .C(net830),
    .X(net139));
 sky130_fd_sc_hd__and2_0 c160 (.A(net128),
    .B(net2),
    .X(net140));
 sky130_fd_sc_hd__and2_0 c161 (.A(net140),
    .B(net134),
    .X(net141));
 sky130_fd_sc_hd__and2_1 c162 (.A(net956),
    .B(net139),
    .X(net142));
 sky130_fd_sc_hd__sdfrbp_1 c163 (.CLK(clknet_leaf_38_clk),
    .D(net131),
    .RESET_B(net137),
    .SCD(net797),
    .SCE(net960),
    .Q(net144),
    .Q_N(net143));
 sky130_fd_sc_hd__sdfbbn_2 c164 (.CLK_N(clknet_leaf_38_clk),
    .D(net137),
    .RESET_B(net142),
    .SCD(net141),
    .SCE(net790),
    .SET_B(net6),
    .Q(net146),
    .Q_N(net145));
 sky130_fd_sc_hd__mux4_2 c165 (.A0(net140),
    .A1(net139),
    .A2(net791),
    .A3(net145),
    .S0(net2),
    .S1(net12),
    .X(net147));
 sky130_fd_sc_hd__edfxbp_1 c166 (.CLK(clknet_leaf_37_clk),
    .D(net147),
    .DE(net11),
    .Q(net149),
    .Q_N(net148));
 sky130_fd_sc_hd__dfbbp_1 c167 (.CLK(clknet_leaf_38_clk),
    .D(net141),
    .RESET_B(net958),
    .SET_B(net139),
    .Q(net151),
    .Q_N(net150));
 sky130_fd_sc_hd__clkbuf_2 c168 (.A(net124),
    .X(net152));
 sky130_fd_sc_hd__and3_1 c169 (.A(net791),
    .B(net793),
    .C(net12),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 c170 (.X(net154));
 sky130_fd_sc_hd__and2_1 c171 (.A(net28),
    .B(net22),
    .X(net155));
 sky130_fd_sc_hd__buf_1 c172 (.A(net725),
    .X(net156));
 sky130_fd_sc_hd__edfxtp_1 c173 (.CLK(clknet_leaf_36_clk),
    .D(net2),
    .DE(net152),
    .Q(net157));
 sky130_fd_sc_hd__sdlclkp_1 c174 (.CLK(clknet_leaf_33_clk),
    .GATE(net111),
    .SCE(net908),
    .GCLK(net158));
 sky130_fd_sc_hd__sdlclkp_2 c175 (.CLK(clknet_leaf_32_clk),
    .GATE(net153),
    .SCE(net888),
    .GCLK(net159));
 sky130_fd_sc_hd__sdlclkp_4 c176 (.CLK(clknet_leaf_39_clk),
    .GATE(net123),
    .SCE(net36),
    .GCLK(net160));
 sky130_fd_sc_hd__or4bb_1 c177 (.A(clknet_1_1__leaf_net158),
    .B(net136),
    .C_N(clknet_1_0__leaf_net160),
    .D_N(net156),
    .X(net161));
 sky130_fd_sc_hd__and2_0 c178 (.A(net136),
    .B(net130),
    .X(net162));
 sky130_fd_sc_hd__dfrbp_1 c179 (.CLK(clknet_leaf_31_clk),
    .D(net155),
    .RESET_B(net156),
    .Q(net164),
    .Q_N(net163));
 sky130_fd_sc_hd__and2_0 c180 (.A(net161),
    .B(clknet_1_0__leaf_net160),
    .X(net165));
 sky130_fd_sc_hd__and2_0 c181 (.A(clknet_1_1__leaf_net158),
    .B(clknet_1_0__leaf_net165),
    .X(net166));
 sky130_fd_sc_hd__and3_1 c182 (.A(net130),
    .B(net25),
    .C(net133),
    .X(net167));
 sky130_fd_sc_hd__mux4_1 c183 (.A0(net167),
    .A1(clknet_1_0__leaf_net158),
    .A2(net157),
    .A3(clknet_1_0__leaf_net166),
    .S0(net36),
    .S1(clknet_1_0__leaf_net165),
    .X(net168));
 sky130_fd_sc_hd__and2_2 c184 (.A(net157),
    .B(net25),
    .X(net169));
 sky130_fd_sc_hd__sdfxbp_1 c185 (.CLK(clknet_leaf_33_clk),
    .D(net167),
    .SCD(clknet_1_0__leaf_net158),
    .SCE(net169),
    .Q(net170));
 sky130_fd_sc_hd__mux4_1 c186 (.A0(net113),
    .A1(net146),
    .A2(net169),
    .A3(net162),
    .S0(net20),
    .S1(clknet_1_1__leaf_net158),
    .X(net171));
 sky130_fd_sc_hd__sdfxbp_1 c187 (.CLK(clknet_leaf_33_clk),
    .D(net894),
    .SCD(net167),
    .SCE(net155),
    .Q(net172));
 sky130_fd_sc_hd__sdfxtp_1 c188 (.CLK(clknet_leaf_32_clk),
    .D(clknet_1_1__leaf_net160),
    .SCD(clknet_1_0__leaf_net171),
    .SCE(net888),
    .Q(net173));
 sky130_fd_sc_hd__buf_1 c189 (.A(net156),
    .X(net174));
 sky130_fd_sc_hd__buf_6 c190 (.A(net58),
    .X(net175));
 sky130_fd_sc_hd__and2_0 c191 (.A(net0),
    .B(net169),
    .X(net176));
 sky130_fd_sc_hd__dfrbp_1 c192 (.CLK(clknet_leaf_32_clk),
    .D(net126),
    .RESET_B(net874),
    .Q(net178),
    .Q_N(net177));
 sky130_fd_sc_hd__sdfxtp_1 c193 (.CLK(clknet_leaf_31_clk),
    .D(net919),
    .SCD(clknet_1_0__leaf_net171),
    .SCE(net25),
    .Q(net179));
 sky130_fd_sc_hd__dfxbp_1 c194 (.CLK(clknet_leaf_12_clk),
    .D(net6),
    .Q(net181),
    .Q_N(net180));
 sky130_fd_sc_hd__dfxbp_1 c195 (.CLK(clknet_leaf_32_clk),
    .D(net176),
    .Q(net182));
 sky130_fd_sc_hd__and2_0 c196 (.A(net845),
    .B(net177),
    .X(net183));
 sky130_fd_sc_hd__and3_1 c197 (.A(net182),
    .B(net45),
    .C(net129),
    .X(net184));
 sky130_fd_sc_hd__dfxtp_1 c198 (.CLK(clknet_leaf_32_clk),
    .D(net176),
    .Q(net185));
 sky130_fd_sc_hd__and2_0 c199 (.A(net45),
    .B(net169),
    .X(net186));
 sky130_fd_sc_hd__sdfxtp_1 c200 (.CLK(clknet_leaf_31_clk),
    .D(net895),
    .SCD(net919),
    .SCE(net6),
    .Q(net187));
 sky130_fd_sc_hd__buf_1 c201 (.A(net173),
    .X(net188));
 sky130_fd_sc_hd__and2_2 c202 (.A(net851),
    .B(net188),
    .X(net189));
 sky130_fd_sc_hd__dfrtn_1 c203 (.CLK_N(clknet_leaf_30_clk),
    .D(net186),
    .RESET_B(net871),
    .Q(net190));
 sky130_fd_sc_hd__dfrtp_1 c204 (.CLK(clknet_leaf_30_clk),
    .D(clknet_1_1__leaf_net171),
    .RESET_B(net852),
    .Q(net191));
 sky130_fd_sc_hd__and2_1 c205 (.A(net872),
    .B(net189),
    .X(net192));
 sky130_fd_sc_hd__dfrtp_1 c206 (.CLK(clknet_leaf_30_clk),
    .D(net186),
    .RESET_B(net190),
    .Q(net193));
 sky130_fd_sc_hd__and2_1 c207 (.A(net189),
    .B(net876),
    .X(net194));
 sky130_fd_sc_hd__dfrtp_1 c208 (.CLK(clknet_leaf_30_clk),
    .D(net106),
    .RESET_B(net194),
    .Q(net195));
 sky130_fd_sc_hd__dfbbn_1 c209 (.CLK_N(clknet_leaf_31_clk),
    .D(net194),
    .RESET_B(net13),
    .SET_B(net174),
    .Q(net197),
    .Q_N(net196));
 sky130_fd_sc_hd__and2_1 c210 (.A(net955),
    .B(net85),
    .X(net198));
 sky130_fd_sc_hd__dfsbp_1 c211 (.CLK(clknet_leaf_27_clk),
    .D(net77),
    .SET_B(net856),
    .Q(net199));
 sky130_fd_sc_hd__and2_0 c212 (.A(net977),
    .B(net83),
    .X(net200));
 sky130_fd_sc_hd__dfsbp_1 c213 (.CLK(clknet_leaf_27_clk),
    .D(net72),
    .SET_B(net860),
    .Q(net202),
    .Q_N(net201));
 sky130_fd_sc_hd__and2_1 c214 (.A(net61),
    .B(net67),
    .X(net203));
 sky130_fd_sc_hd__and2_0 c215 (.A(net110),
    .B(net83),
    .X(net204));
 sky130_fd_sc_hd__dfstp_1 c216 (.CLK(clknet_leaf_30_clk),
    .D(net198),
    .SET_B(net864),
    .Q(net205));
 sky130_fd_sc_hd__dfstp_1 c217 (.CLK(clknet_leaf_21_clk),
    .D(net902),
    .SET_B(net135),
    .Q(net206));
 sky130_fd_sc_hd__dfstp_1 c218 (.CLK(clknet_leaf_29_clk),
    .D(net192),
    .SET_B(net858),
    .Q(net207));
 sky130_fd_sc_hd__and2_0 c219 (.A(net195),
    .B(net60),
    .X(net208));
 sky130_fd_sc_hd__and2_1 c220 (.A(net200),
    .B(net203),
    .X(net209));
 sky130_fd_sc_hd__dlrbn_1 c221 (.D(net64),
    .GATE_N(clknet_leaf_30_clk),
    .RESET_B(net192),
    .Q(net211),
    .Q_N(net210));
 sky130_fd_sc_hd__and2_1 c222 (.A(net208),
    .B(net200),
    .X(net212));
 sky130_fd_sc_hd__and2_1 c223 (.A(net207),
    .B(net204),
    .X(net213));
 sky130_fd_sc_hd__dlrbn_1 c224 (.D(net947),
    .GATE_N(clknet_leaf_27_clk),
    .RESET_B(net209),
    .Q(net215),
    .Q_N(net214));
 sky130_fd_sc_hd__dlrbp_2 c225 (.D(net36),
    .GATE(clknet_leaf_30_clk),
    .RESET_B(net152),
    .Q(net820),
    .Q_N(net216));
 sky130_fd_sc_hd__and2_0 c226 (.A(net204),
    .B(net818),
    .X(net217));
 sky130_fd_sc_hd__dfbbn_1 c227 (.CLK_N(clknet_leaf_30_clk),
    .D(net152),
    .RESET_B(net879),
    .SET_B(net216),
    .Q(net218));
 sky130_fd_sc_hd__dlrbp_1 c228 (.D(net991),
    .GATE(clknet_leaf_21_clk),
    .RESET_B(net198),
    .Q(net220),
    .Q_N(net219));
 sky130_fd_sc_hd__dfbbp_1 c229 (.CLK(clknet_leaf_27_clk),
    .D(net217),
    .RESET_B(net4),
    .SET_B(net861),
    .Q(net221));
 sky130_fd_sc_hd__a2111o_1 c230 (.A1(net221),
    .A2(net212),
    .B1(net216),
    .C1(net189),
    .D1(net203),
    .X(net222));
 sky130_fd_sc_hd__sdfxbp_1 c231 (.CLK(clknet_leaf_27_clk),
    .D(net786),
    .SCD(net213),
    .SCE(net966),
    .Q(net223));
 sky130_fd_sc_hd__dlrtn_1 c232 (.D(net105),
    .GATE_N(clknet_leaf_27_clk),
    .RESET_B(net916),
    .Q(net224));
 sky130_fd_sc_hd__and2_0 c233 (.A(net223),
    .B(net88),
    .X(net225));
 sky130_fd_sc_hd__and2_0 c234 (.A(net85),
    .B(net203),
    .X(net226));
 sky130_fd_sc_hd__dlrtn_1 c235 (.D(net209),
    .GATE_N(clknet_leaf_26_clk),
    .RESET_B(net224),
    .Q(net812));
 sky130_fd_sc_hd__dlrtn_1 c236 (.D(net213),
    .GATE_N(clknet_leaf_27_clk),
    .RESET_B(net978),
    .Q(net227));
 sky130_fd_sc_hd__sdfxbp_1 c237 (.CLK(clknet_leaf_28_clk),
    .D(net903),
    .SCD(net105),
    .SCE(net995),
    .Q(net228));
 sky130_fd_sc_hd__and2_1 c238 (.A(net104),
    .B(net789),
    .X(net229));
 sky130_fd_sc_hd__dlrtp_1 c239 (.D(net226),
    .GATE(clknet_leaf_26_clk),
    .RESET_B(net209),
    .Q(net230));
 sky130_fd_sc_hd__or4bb_1 c240 (.A(net225),
    .B(net85),
    .C_N(net230),
    .D_N(net229),
    .X(net231));
 sky130_fd_sc_hd__dlrtp_1 c241 (.D(net231),
    .GATE(clknet_leaf_26_clk),
    .RESET_B(net230),
    .Q(net232));
 sky130_fd_sc_hd__and3_1 c242 (.A(net227),
    .B(net205),
    .C(net786),
    .X(net233));
 sky130_fd_sc_hd__dlrtp_1 c243 (.D(net83),
    .GATE(clknet_leaf_26_clk),
    .RESET_B(net231),
    .Q(net234));
 sky130_fd_sc_hd__and3_1 c244 (.A(net968),
    .B(net230),
    .C(net229),
    .X(net235));
 sky130_fd_sc_hd__and2_0 c245 (.A(net203),
    .B(net973),
    .X(net236));
 sky130_fd_sc_hd__and2_0 c246 (.A(net75),
    .B(net234),
    .X(net237));
 sky130_fd_sc_hd__edfxbp_1 c247 (.CLK(clknet_leaf_26_clk),
    .D(net236),
    .DE(net104),
    .Q(net238));
 sky130_fd_sc_hd__or4bb_1 c248 (.A(net237),
    .B(net55),
    .C_N(net229),
    .D_N(net85),
    .X(net239));
 sky130_fd_sc_hd__edfxtp_1 c249 (.CLK(clknet_leaf_26_clk),
    .D(net239),
    .DE(net831),
    .Q(net240));
 sky130_fd_sc_hd__and2_0 c25 (.A(net799),
    .B(net801),
    .X(net0));
 sky130_fd_sc_hd__mux4_1 c250 (.A0(net233),
    .A1(net813),
    .A2(net99),
    .A3(net229),
    .S0(net240),
    .S1(net237),
    .X(net241));
 sky130_fd_sc_hd__sdlclkp_1 c251 (.CLK(clknet_leaf_25_clk),
    .GATE(net235),
    .SCE(net239),
    .GCLK(net242));
 sky130_fd_sc_hd__buf_1 c252 (.A(net807),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_1 c253 (.A(net122),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_1 c254 (.A(net122),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_1 c255 (.A(net922),
    .X(net246));
 sky130_fd_sc_hd__dlymetal6s2s_1 c256 (.A(net244),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_1 c257 (.A(net245),
    .X(net248));
 sky130_fd_sc_hd__and2_4 c258 (.A(net785),
    .B(net247),
    .X(net249));
 sky130_fd_sc_hd__sdlclkp_2 c259 (.CLK(clknet_leaf_3_clk),
    .GATE(net109),
    .SCE(net126),
    .GCLK(net250));
 sky130_fd_sc_hd__and2_2 c26 (.A(net805),
    .B(net803),
    .X(net1));
 sky130_fd_sc_hd__and2_0 c260 (.A(net808),
    .B(clknet_1_0__leaf_net250),
    .X(net251));
 sky130_fd_sc_hd__buf_1 c261 (.A(clknet_1_1__leaf_net250),
    .X(net252));
 sky130_fd_sc_hd__and2_0 c262 (.A(clknet_1_0__leaf_net252),
    .B(clknet_1_1__leaf_net251),
    .X(net253));
 sky130_fd_sc_hd__buf_1 c263 (.A(net797),
    .X(net254));
 sky130_fd_sc_hd__buf_1 c264 (.A(clknet_1_0__leaf_net253),
    .X(net255));
 sky130_fd_sc_hd__buf_1 c265 (.A(net254),
    .X(net256));
 sky130_fd_sc_hd__and2_1 c266 (.A(net256),
    .B(net254),
    .X(net257));
 sky130_fd_sc_hd__and3_1 c267 (.A(net248),
    .B(clknet_1_0__leaf_net250),
    .C(net244),
    .X(net258));
 sky130_fd_sc_hd__buf_1 c268 (.A(net254),
    .X(net259));
 sky130_fd_sc_hd__and3_1 c269 (.A(net243),
    .B(net259),
    .C(clknet_1_1__leaf_net251),
    .X(net260));
 sky130_fd_sc_hd__and2_1 c27 (.A(net801),
    .B(net798),
    .X(net2));
 sky130_fd_sc_hd__sdlclkp_4 c270 (.CLK(clknet_leaf_3_clk),
    .GATE(clknet_1_0__leaf_net260),
    .SCE(net787),
    .GCLK(net261));
 sky130_fd_sc_hd__buf_2 c271 (.A(net922),
    .X(net262));
 sky130_fd_sc_hd__mux4_1 c272 (.A0(clknet_1_1__leaf_net258),
    .A1(clknet_1_0__leaf_net261),
    .A2(net108),
    .A3(clknet_1_1__leaf_net251),
    .S0(net262),
    .S1(net256),
    .X(net263));
 sky130_fd_sc_hd__and2_1 c273 (.A(net11),
    .B(net909),
    .X(net264));
 sky130_fd_sc_hd__buf_1 c274 (.A(net16),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_1 c275 (.A(net751),
    .X(net266));
 sky130_fd_sc_hd__and2_2 c276 (.A(net151),
    .B(net259),
    .X(net267));
 sky130_fd_sc_hd__buf_2 c277 (.A(net751),
    .X(net829));
 sky130_fd_sc_hd__dfrbp_1 c278 (.CLK(clknet_leaf_6_clk),
    .D(net142),
    .RESET_B(net147),
    .Q(net269),
    .Q_N(net268));
 sky130_fd_sc_hd__and2_2 c279 (.A(net264),
    .B(net834),
    .X(net270));
 sky130_fd_sc_hd__and2_1 c28 (.A(net0),
    .B(net804),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 c280 (.A(net920),
    .X(net271));
 sky130_fd_sc_hd__dfrbp_1 c281 (.CLK(clknet_leaf_37_clk),
    .D(net270),
    .RESET_B(net15),
    .Q(net273),
    .Q_N(net272));
 sky130_fd_sc_hd__and2_1 c282 (.A(net245),
    .B(net247),
    .X(net274));
 sky130_fd_sc_hd__dfrtn_1 c283 (.CLK_N(clknet_leaf_37_clk),
    .D(net797),
    .RESET_B(net257),
    .Q(net275));
 sky130_fd_sc_hd__and2_1 c284 (.A(net139),
    .B(net264),
    .X(net276));
 sky130_fd_sc_hd__and2_0 c285 (.A(net982),
    .B(net275),
    .X(net277));
 sky130_fd_sc_hd__and2_0 c286 (.A(net846),
    .B(net275),
    .X(net278));
 sky130_fd_sc_hd__sdfxtp_1 c287 (.CLK(clknet_leaf_37_clk),
    .D(net278),
    .SCD(net275),
    .SCE(net834),
    .Q(net279));
 sky130_fd_sc_hd__mux4_1 c288 (.A0(net279),
    .A1(net148),
    .A2(net272),
    .A3(net277),
    .S0(net270),
    .S1(net834),
    .X(net280));
 sky130_fd_sc_hd__sdfxtp_2 c289 (.CLK(clknet_leaf_37_clk),
    .D(net277),
    .SCD(net267),
    .SCE(net760),
    .Q(net281));
 sky130_fd_sc_hd__and2_2 c29 (.A(net800),
    .B(net799),
    .X(net818));
 sky130_fd_sc_hd__dfrtp_1 c290 (.CLK(clknet_leaf_37_clk),
    .D(net271),
    .RESET_B(net278),
    .Q(net282));
 sky130_fd_sc_hd__dfrtp_1 c291 (.CLK(clknet_leaf_37_clk),
    .D(net907),
    .RESET_B(net127),
    .Q(net283));
 sky130_fd_sc_hd__and3_2 c292 (.A(net279),
    .B(net283),
    .C(net761),
    .X(net284));
 sky130_fd_sc_hd__and3_2 c293 (.A(net265),
    .B(net907),
    .C(net921),
    .X(net285));
 sky130_fd_sc_hd__and2_1 c294 (.A(net162),
    .B(net146),
    .X(net286));
 sky130_fd_sc_hd__and3_1 c295 (.A(net13),
    .B(net110),
    .C(clknet_1_1__leaf_net250),
    .X(net287));
 sky130_fd_sc_hd__sdfbbn_1 c296 (.CLK_N(clknet_leaf_39_clk),
    .D(net155),
    .RESET_B(net990),
    .SCD(clknet_1_0__leaf_net251),
    .SCE(net274),
    .SET_B(net834),
    .Q(net288));
 sky130_fd_sc_hd__and2_1 c297 (.A(net286),
    .B(net22),
    .X(net289));
 sky130_fd_sc_hd__and2_0 c298 (.A(clknet_1_0__leaf_net251),
    .B(net285),
    .X(net290));
 sky130_fd_sc_hd__buf_1 c299 (.A(net743),
    .X(net291));
 sky130_fd_sc_hd__and2_2 c30 (.A(net818),
    .B(net805),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 c300 (.A(net743),
    .X(net292));
 sky130_fd_sc_hd__dfrtp_4 c301 (.CLK(clknet_leaf_39_clk),
    .D(net921),
    .RESET_B(clknet_1_0__leaf_net290),
    .Q(net293));
 sky130_fd_sc_hd__and2_2 c302 (.A(net803),
    .B(net292),
    .X(net828));
 sky130_fd_sc_hd__a2111o_1 c303 (.A1(net790),
    .A2(net286),
    .B1(net791),
    .C1(net22),
    .D1(clknet_1_0__leaf_net165),
    .X(net294));
 sky130_fd_sc_hd__mux4_1 c304 (.A0(clknet_1_1__leaf_net290),
    .A1(clknet_1_0__leaf_net294),
    .A2(net291),
    .A3(net293),
    .S0(net147),
    .S1(net270),
    .X(net295));
 sky130_fd_sc_hd__sdfxtp_2 c305 (.CLK(clknet_leaf_39_clk),
    .D(net275),
    .SCD(net162),
    .SCE(clknet_1_0__leaf_net290),
    .Q(net296));
 sky130_fd_sc_hd__and2_0 c306 (.A(net159),
    .B(net296),
    .X(net297));
 sky130_fd_sc_hd__and2_2 c307 (.A(net172),
    .B(net296),
    .X(net298));
 sky130_fd_sc_hd__and3_1 c308 (.A(net22),
    .B(net293),
    .C(net282),
    .X(net299));
 sky130_fd_sc_hd__and2_2 c309 (.A(net288),
    .B(net129),
    .X(net811));
 sky130_fd_sc_hd__and2_4 c31 (.A(net801),
    .B(net0),
    .X(net5));
 sky130_fd_sc_hd__dfbbn_1 c310 (.CLK_N(clknet_leaf_0_clk),
    .D(net20),
    .RESET_B(net249),
    .SET_B(net298),
    .Q(net301),
    .Q_N(net300));
 sky130_fd_sc_hd__dfbbn_1 c311 (.CLK_N(clknet_leaf_0_clk),
    .D(clknet_1_0__leaf_net294),
    .RESET_B(net912),
    .SET_B(net293),
    .Q(net302));
 sky130_fd_sc_hd__and2_1 c312 (.A(net302),
    .B(net286),
    .X(net303));
 sky130_fd_sc_hd__a2111o_1 c313 (.A1(net298),
    .A2(net20),
    .B1(net300),
    .C1(clknet_1_0__leaf_net165),
    .D1(net291),
    .X(net304));
 sky130_fd_sc_hd__dfsbp_1 c314 (.CLK(clknet_leaf_32_clk),
    .D(net267),
    .SET_B(net762),
    .Q(net306),
    .Q_N(net305));
 sky130_fd_sc_hd__mux4_1 c315 (.A0(net174),
    .A1(net49),
    .A2(net184),
    .A3(net285),
    .S0(net298),
    .S1(net169),
    .X(net307));
 sky130_fd_sc_hd__and2_0 c316 (.A(net979),
    .B(net756),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_1 c317 (.A(net745),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_1 c318 (.A(net744),
    .X(net310));
 sky130_fd_sc_hd__and2_0 c319 (.A(net129),
    .B(net25),
    .X(net311));
 sky130_fd_sc_hd__and2_2 c32 (.A(net3),
    .B(net4),
    .X(net6));
 sky130_fd_sc_hd__and2_0 c320 (.A(net188),
    .B(net828),
    .X(net312));
 sky130_fd_sc_hd__and2_1 c321 (.A(net291),
    .B(net945),
    .X(net313));
 sky130_fd_sc_hd__dfsbp_1 c322 (.CLK(clknet_leaf_30_clk),
    .D(clknet_1_1__leaf_net294),
    .SET_B(net285),
    .Q(net314));
 sky130_fd_sc_hd__and2_0 c323 (.A(net169),
    .B(net183),
    .X(net315));
 sky130_fd_sc_hd__and2_0 c324 (.A(net306),
    .B(net293),
    .X(net316));
 sky130_fd_sc_hd__and2_1 c325 (.A(net183),
    .B(net311),
    .X(net317));
 sky130_fd_sc_hd__dfbbp_1 c326 (.CLK(clknet_leaf_20_clk),
    .D(net890),
    .RESET_B(net317),
    .SET_B(clknet_1_1__leaf_net294),
    .Q(net319),
    .Q_N(net318));
 sky130_fd_sc_hd__sdfxbp_1 c327 (.CLK(clknet_leaf_31_clk),
    .D(net317),
    .SCD(net49),
    .SCE(net188),
    .Q(net321),
    .Q_N(net320));
 sky130_fd_sc_hd__and2_0 c328 (.A(net314),
    .B(net298),
    .X(net322));
 sky130_fd_sc_hd__dfstp_1 c329 (.CLK(clknet_leaf_31_clk),
    .D(net980),
    .SET_B(net317),
    .Q(net323));
 sky130_fd_sc_hd__buf_1 c33 (.A(net790),
    .X(net7));
 sky130_fd_sc_hd__and2_2 c330 (.A(net875),
    .B(net189),
    .X(net324));
 sky130_fd_sc_hd__sdfrtn_1 c331 (.CLK_N(clknet_leaf_21_clk),
    .D(net319),
    .RESET_B(net191),
    .SCD(net324),
    .SCE(net317),
    .Q(net325));
 sky130_fd_sc_hd__dfstp_1 c332 (.CLK(clknet_leaf_21_clk),
    .D(net325),
    .SET_B(net324),
    .Q(net326));
 sky130_fd_sc_hd__and2_0 c333 (.A(net322),
    .B(net169),
    .X(net327));
 sky130_fd_sc_hd__mux4_1 c334 (.A0(net316),
    .A1(net320),
    .A2(net315),
    .A3(net326),
    .S0(net291),
    .S1(net121),
    .X(net328));
 sky130_fd_sc_hd__and2_2 c335 (.A(net311),
    .B(net756),
    .X(net833));
 sky130_fd_sc_hd__and2_1 c336 (.A(net281),
    .B(net764),
    .X(net329));
 sky130_fd_sc_hd__and2_0 c337 (.A(net312),
    .B(net329),
    .X(net330));
 sky130_fd_sc_hd__buf_1 c338 (.A(net899),
    .X(net331));
 sky130_fd_sc_hd__and2_0 c339 (.A(net298),
    .B(net923),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_4 c34 (.A(net1),
    .X(net8));
 sky130_fd_sc_hd__sdfxbp_1 c340 (.CLK(clknet_leaf_23_clk),
    .D(net913),
    .SCD(net834),
    .SCE(net831),
    .Q(net333));
 sky130_fd_sc_hd__clkbuf_1 c341 (.A(net747),
    .X(net334));
 sky130_fd_sc_hd__and3_1 c342 (.A(net191),
    .B(net329),
    .C(net219),
    .X(net335));
 sky130_fd_sc_hd__and3_1 c343 (.A(net971),
    .B(net820),
    .C(net803),
    .X(net336));
 sky130_fd_sc_hd__sdfxtp_1 c344 (.CLK(clknet_leaf_21_clk),
    .D(net222),
    .SCD(net913),
    .SCE(net907),
    .Q(net337));
 sky130_fd_sc_hd__sdfxtp_1 c345 (.CLK(clknet_leaf_21_clk),
    .D(net135),
    .SCD(net329),
    .SCE(net222),
    .Q(net338));
 sky130_fd_sc_hd__and2_0 c346 (.A(net334),
    .B(net220),
    .X(net339));
 sky130_fd_sc_hd__dfstp_1 c347 (.CLK(clknet_leaf_21_clk),
    .D(net313),
    .SET_B(net135),
    .Q(net340));
 sky130_fd_sc_hd__and2_0 c348 (.A(net333),
    .B(net340),
    .X(net341));
 sky130_fd_sc_hd__sdfxtp_1 c349 (.CLK(clknet_leaf_21_clk),
    .D(net336),
    .SCD(net943),
    .SCE(net82),
    .Q(net342));
 sky130_fd_sc_hd__and3_1 c35 (.A(net798),
    .B(net1),
    .C(net8),
    .X(net9));
 sky130_fd_sc_hd__and2_1 c350 (.A(net341),
    .B(net828),
    .X(net343));
 sky130_fd_sc_hd__and3_1 c351 (.A(net881),
    .B(net67),
    .C(net340),
    .X(net344));
 sky130_fd_sc_hd__or4bb_4 c352 (.A(net332),
    .B(net834),
    .C_N(net343),
    .D_N(net189),
    .X(net345));
 sky130_fd_sc_hd__dfbbn_1 c353 (.CLK_N(clknet_leaf_21_clk),
    .D(net833),
    .RESET_B(net340),
    .SET_B(net763),
    .Q(net347),
    .Q_N(net346));
 sky130_fd_sc_hd__dfbbn_1 c354 (.CLK_N(clknet_leaf_21_clk),
    .D(net25),
    .RESET_B(net189),
    .SET_B(net345),
    .Q(net349),
    .Q_N(net348));
 sky130_fd_sc_hd__and2_0 c355 (.A(net339),
    .B(net953),
    .X(net350));
 sky130_fd_sc_hd__dfbbp_1 c356 (.CLK(clknet_leaf_22_clk),
    .D(net82),
    .RESET_B(net346),
    .SET_B(net345),
    .Q(net352),
    .Q_N(net351));
 sky130_fd_sc_hd__and2_1 c357 (.A(net212),
    .B(net826),
    .X(net809));
 sky130_fd_sc_hd__dlrbn_1 c358 (.D(net289),
    .GATE_N(clknet_leaf_23_clk),
    .RESET_B(net850),
    .Q(net353));
 sky130_fd_sc_hd__and2_0 c359 (.A(net5),
    .B(net758),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_2 c36 (.A(net732),
    .X(net10));
 sky130_fd_sc_hd__dlrbn_1 c360 (.D(net232),
    .GATE_N(clknet_leaf_25_clk),
    .RESET_B(net831),
    .Q(net355));
 sky130_fd_sc_hd__and2_0 c361 (.A(net297),
    .B(clknet_1_1__leaf_net242),
    .X(net356));
 sky130_fd_sc_hd__dlrbp_1 c362 (.D(net98),
    .GATE(clknet_leaf_25_clk),
    .RESET_B(net232),
    .Q(net358),
    .Q_N(net357));
 sky130_fd_sc_hd__and3_1 c363 (.A(net95),
    .B(net810),
    .C(clknet_1_0__leaf_net356),
    .X(net359));
 sky130_fd_sc_hd__sdfxbp_1 c364 (.CLK(clknet_leaf_24_clk),
    .D(clknet_1_0__leaf_net359),
    .SCD(net918),
    .SCE(net99),
    .Q(net361),
    .Q_N(net360));
 sky130_fd_sc_hd__and2_0 c365 (.A(net932),
    .B(net212),
    .X(net362));
 sky130_fd_sc_hd__and3_1 c366 (.A(net229),
    .B(net358),
    .C(net360),
    .X(net363));
 sky130_fd_sc_hd__dlrbp_1 c367 (.D(net99),
    .GATE(clknet_leaf_24_clk),
    .RESET_B(net8),
    .Q(net364));
 sky130_fd_sc_hd__dlrtn_1 c368 (.D(net353),
    .GATE_N(clknet_leaf_23_clk),
    .RESET_B(net809),
    .Q(net365));
 sky130_fd_sc_hd__and3_1 c369 (.A(net365),
    .B(net364),
    .C(net338),
    .X(net366));
 sky130_fd_sc_hd__and2_1 c37 (.A(net806),
    .B(net10),
    .X(net11));
 sky130_fd_sc_hd__sdfxbp_1 c370 (.CLK(clknet_leaf_23_clk),
    .D(net350),
    .SCD(net957),
    .SCE(net345),
    .Q(net367));
 sky130_fd_sc_hd__and3_1 c371 (.A(net986),
    .B(net229),
    .C(net365),
    .X(net368));
 sky130_fd_sc_hd__and3_1 c372 (.A(net285),
    .B(net361),
    .C(net366),
    .X(net369));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net369),
    .A1(net354),
    .A2(net345),
    .A3(net365),
    .S0(net358),
    .S1(clknet_1_1__leaf_net356),
    .X(net370));
 sky130_fd_sc_hd__sdfxtp_1 c374 (.CLK(clknet_leaf_23_clk),
    .D(net368),
    .SCD(net343),
    .SCE(net972),
    .Q(net371));
 sky130_fd_sc_hd__sdfxtp_1 c375 (.CLK(clknet_leaf_24_clk),
    .D(net918),
    .SCD(clknet_1_0__leaf_net359),
    .SCE(net765),
    .Q(net372));
 sky130_fd_sc_hd__mux4_1 c376 (.A0(net345),
    .A1(net363),
    .A2(clknet_1_1__leaf_net359),
    .A3(net788),
    .S0(net357),
    .S1(net365),
    .X(net373));
 sky130_fd_sc_hd__mux4_1 c377 (.A0(net367),
    .A1(net371),
    .A2(net365),
    .A3(clknet_1_1__leaf_net359),
    .S0(net357),
    .S1(net363),
    .X(net374));
 sky130_fd_sc_hd__and2_2 c378 (.A(net119),
    .B(net120),
    .X(net375));
 sky130_fd_sc_hd__dlymetal6s2s_1 c379 (.A(net738),
    .X(net376));
 sky130_fd_sc_hd__and3_4 c38 (.A(net11),
    .B(net1),
    .C(net7),
    .X(net12));
 sky130_fd_sc_hd__buf_1 c380 (.A(net244),
    .X(net377));
 sky130_fd_sc_hd__dlymetal6s2s_1 c381 (.A(net739),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_4 c382 (.A(net378),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_4 c383 (.A(net846),
    .X(net380));
 sky130_fd_sc_hd__buf_2 c384 (.A(net375),
    .X(net381));
 sky130_fd_sc_hd__and2_1 c385 (.A(net381),
    .B(net379),
    .X(net382));
 sky130_fd_sc_hd__dlrtn_1 c386 (.D(net257),
    .GATE_N(clknet_leaf_3_clk),
    .RESET_B(net382),
    .Q(net383));
 sky130_fd_sc_hd__dlrtn_1 c387 (.D(net376),
    .GATE_N(clknet_leaf_1_clk),
    .RESET_B(clknet_1_0__leaf_net255),
    .Q(net384));
 sky130_fd_sc_hd__dlrtp_2 c388 (.D(net382),
    .GATE(clknet_leaf_4_clk),
    .RESET_B(net381),
    .Q(net385));
 sky130_fd_sc_hd__buf_1 c389 (.A(net379),
    .X(net386));
 sky130_fd_sc_hd__dlymetal6s2s_1 c39 (.A(net731),
    .X(net13));
 sky130_fd_sc_hd__and2_1 c390 (.A(net384),
    .B(net379),
    .X(net387));
 sky130_fd_sc_hd__mux4_1 c391 (.A0(net386),
    .A1(net387),
    .A2(net377),
    .A3(clknet_1_1__leaf_net255),
    .S0(net380),
    .S1(net379),
    .X(net388));
 sky130_fd_sc_hd__and2_1 c392 (.A(net248),
    .B(net768),
    .X(net389));
 sky130_fd_sc_hd__and2_0 c393 (.A(net376),
    .B(net759),
    .X(net390));
 sky130_fd_sc_hd__and2_0 c394 (.A(net950),
    .B(net381),
    .X(net391));
 sky130_fd_sc_hd__dlrtp_1 c395 (.D(net389),
    .GATE(clknet_leaf_4_clk),
    .RESET_B(net391),
    .Q(net392));
 sky130_fd_sc_hd__dlrtp_2 c396 (.D(net391),
    .GATE(clknet_leaf_3_clk),
    .RESET_B(net392),
    .Q(net393));
 sky130_fd_sc_hd__sdfxtp_1 c397 (.CLK(clknet_leaf_3_clk),
    .D(net389),
    .SCD(net963),
    .SCE(net931),
    .Q(net394));
 sky130_fd_sc_hd__dfbbn_1 c398 (.CLK_N(clknet_leaf_3_clk),
    .D(clknet_1_0__leaf_net390),
    .RESET_B(net394),
    .SET_B(net389),
    .Q(net396),
    .Q_N(net395));
 sky130_fd_sc_hd__clkbuf_1 c399 (.A(net737),
    .X(net397));
 sky130_fd_sc_hd__and3_2 c40 (.A(net12),
    .B(net798),
    .C(net803),
    .X(net14));
 sky130_fd_sc_hd__and2_0 c400 (.A(net266),
    .B(clknet_1_0__leaf_net261),
    .X(net398));
 sky130_fd_sc_hd__and2_0 c401 (.A(clknet_1_1__leaf_net261),
    .B(net800),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_1 c402 (.A(net737),
    .X(net400));
 sky130_fd_sc_hd__and3_1 c403 (.A(clknet_1_1__leaf_net398),
    .B(net5),
    .C(net397),
    .X(net401));
 sky130_fd_sc_hd__and3_1 c404 (.A(clknet_1_1__leaf_net399),
    .B(net138),
    .C(net393),
    .X(net402));
 sky130_fd_sc_hd__and2_2 c405 (.A(net259),
    .B(net115),
    .X(net403));
 sky130_fd_sc_hd__edfxbp_1 c406 (.CLK(clknet_leaf_1_clk),
    .D(net246),
    .DE(net276),
    .Q(net405),
    .Q_N(net404));
 sky130_fd_sc_hd__dfbbn_1 c407 (.CLK_N(clknet_leaf_3_clk),
    .D(net256),
    .RESET_B(net396),
    .SET_B(clknet_1_0__leaf_net402),
    .Q(net407),
    .Q_N(net406));
 sky130_fd_sc_hd__edfxtp_1 c408 (.CLK(clknet_leaf_1_clk),
    .D(net397),
    .DE(net403),
    .Q(net408));
 sky130_fd_sc_hd__dfbbp_1 c409 (.CLK(clknet_leaf_1_clk),
    .D(clknet_1_0__leaf_net402),
    .RESET_B(net395),
    .SET_B(net936),
    .Q(net410),
    .Q_N(net409));
 sky130_fd_sc_hd__dfbbn_1 c41 (.CLK_N(clknet_leaf_36_clk),
    .D(net14),
    .RESET_B(net12),
    .SET_B(net3),
    .Q(net16),
    .Q_N(net15));
 sky130_fd_sc_hd__and2_0 c410 (.A(net119),
    .B(net116),
    .X(net411));
 sky130_fd_sc_hd__and2_2 c411 (.A(net411),
    .B(net404),
    .X(net412));
 sky130_fd_sc_hd__and3_1 c412 (.A(clknet_1_0__leaf_net399),
    .B(net409),
    .C(net412),
    .X(net413));
 sky130_fd_sc_hd__and2_0 c413 (.A(net412),
    .B(net408),
    .X(net414));
 sky130_fd_sc_hd__sdfxbp_1 c414 (.CLK(clknet_leaf_4_clk),
    .D(net790),
    .SCD(net877),
    .SCE(net403),
    .Q(net415));
 sky130_fd_sc_hd__sdfxbp_1 c415 (.CLK(clknet_leaf_1_clk),
    .D(net414),
    .SCD(net412),
    .SCE(net883),
    .Q(net416));
 sky130_fd_sc_hd__and2_0 c416 (.A(net410),
    .B(net411),
    .X(net417));
 sky130_fd_sc_hd__sdfbbp_1 c417 (.CLK(clknet_leaf_1_clk),
    .D(net901),
    .RESET_B(net417),
    .SCD(net400),
    .SCE(net403),
    .SET_B(clknet_1_0__leaf_net398),
    .Q(net418));
 sky130_fd_sc_hd__sdfbbn_1 c418 (.CLK_N(clknet_leaf_1_clk),
    .D(net418),
    .RESET_B(clknet_1_1__leaf_net402),
    .SCD(net385),
    .SCE(net375),
    .SET_B(net380),
    .Q(net420),
    .Q_N(net419));
 sky130_fd_sc_hd__a2111o_1 c419 (.A1(net406),
    .A2(net420),
    .B1(net408),
    .C1(net264),
    .D1(net412),
    .X(net421));
 sky130_fd_sc_hd__buf_1 c42 (.A(net795),
    .X(net17));
 sky130_fd_sc_hd__sdfxtp_1 c420 (.CLK(clknet_leaf_0_clk),
    .D(net304),
    .SCD(net381),
    .SCE(clknet_1_0__leaf_net757),
    .Q(net422));
 sky130_fd_sc_hd__clkbuf_1 c421 (.A(net727),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_1 c422 (.A(net726),
    .X(net424));
 sky130_fd_sc_hd__sdlclkp_1 c423 (.CLK(clknet_leaf_0_clk),
    .GATE(net954),
    .SCE(net274),
    .GCLK(net425));
 sky130_fd_sc_hd__sdlclkp_2 c424 (.CLK(clknet_leaf_0_clk),
    .GATE(clknet_1_0__leaf_net401),
    .SCE(net262),
    .GCLK(net426));
 sky130_fd_sc_hd__sdlclkp_4 c425 (.CLK(clknet_leaf_11_clk),
    .GATE(net126),
    .SCE(net300),
    .GCLK(net427));
 sky130_fd_sc_hd__dfrbp_1 c426 (.CLK(clknet_leaf_19_clk),
    .D(net303),
    .RESET_B(net834),
    .Q(net429),
    .Q_N(net428));
 sky130_fd_sc_hd__sdfxtp_1 c427 (.CLK(clknet_leaf_0_clk),
    .D(net270),
    .SCD(net126),
    .SCE(clknet_1_0__leaf_net757),
    .Q(net430));
 sky130_fd_sc_hd__and2_0 c428 (.A(net423),
    .B(net26),
    .X(net431));
 sky130_fd_sc_hd__and2_0 c429 (.A(net425),
    .B(net143),
    .X(net432));
 sky130_fd_sc_hd__buf_1 c43 (.A(net798),
    .X(net18));
 sky130_fd_sc_hd__dfrbp_1 c430 (.CLK(clknet_leaf_11_clk),
    .D(net407),
    .RESET_B(net126),
    .Q(net434),
    .Q_N(net433));
 sky130_fd_sc_hd__and3_1 c431 (.A(net384),
    .B(net375),
    .C(net429),
    .X(net435));
 sky130_fd_sc_hd__dfrtn_1 c432 (.CLK_N(clknet_leaf_0_clk),
    .D(net400),
    .RESET_B(clknet_1_1__leaf_net166),
    .Q(net436));
 sky130_fd_sc_hd__dfrtp_1 c433 (.CLK(clknet_leaf_1_clk),
    .D(clknet_1_1__leaf_net390),
    .RESET_B(clknet_1_1__leaf_net401),
    .Q(net437));
 sky130_fd_sc_hd__dfrtp_1 c434 (.CLK(clknet_leaf_0_clk),
    .D(clknet_1_0__leaf_net166),
    .RESET_B(clknet_1_0__leaf_net432),
    .Q(net438));
 sky130_fd_sc_hd__sdfxtp_1 c435 (.CLK(clknet_leaf_19_clk),
    .D(net412),
    .SCD(net435),
    .SCE(net249),
    .Q(net439));
 sky130_fd_sc_hd__dfrtp_4 c436 (.CLK(clknet_leaf_0_clk),
    .D(net274),
    .RESET_B(net270),
    .Q(net440));
 sky130_fd_sc_hd__and2_0 c437 (.A(net431),
    .B(net436),
    .X(net441));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(net441),
    .A1(net435),
    .A2(net303),
    .A3(net440),
    .S0(net422),
    .S1(net818),
    .X(net442));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net435),
    .A1(net26),
    .A2(net433),
    .A3(net830),
    .S0(net440),
    .S1(net769),
    .X(net443));
 sky130_fd_sc_hd__buf_1 c44 (.A(net796),
    .X(net19));
 sky130_fd_sc_hd__dfbbn_1 c440 (.CLK_N(clknet_leaf_12_clk),
    .D(net443),
    .RESET_B(net412),
    .SET_B(net770),
    .Q(net444));
 sky130_fd_sc_hd__and3_1 c441 (.A(net434),
    .B(clknet_1_1__leaf_net432),
    .C(net408),
    .X(net445));
 sky130_fd_sc_hd__and2_1 c442 (.A(net197),
    .B(net408),
    .X(net446));
 sky130_fd_sc_hd__and3_1 c443 (.A(net422),
    .B(net309),
    .C(clknet_1_0__leaf_net287),
    .X(net447));
 sky130_fd_sc_hd__and2_0 c444 (.A(net437),
    .B(net318),
    .X(net448));
 sky130_fd_sc_hd__and2_0 c445 (.A(net326),
    .B(clknet_1_1__leaf_net287),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_1 c446 (.A(net741),
    .X(net450));
 sky130_fd_sc_hd__dfbbn_1 c447 (.CLK_N(clknet_leaf_20_clk),
    .D(net426),
    .RESET_B(net324),
    .SET_B(net927),
    .Q(net452),
    .Q_N(net451));
 sky130_fd_sc_hd__dfbbp_1 c448 (.CLK(clknet_leaf_20_clk),
    .D(net49),
    .RESET_B(net326),
    .SET_B(net249),
    .Q(net454),
    .Q_N(net453));
 sky130_fd_sc_hd__clkbuf_1 c449 (.A(net742),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_2 c45 (.A(net19),
    .X(net20));
 sky130_fd_sc_hd__sdfbbn_1 c450 (.CLK_N(clknet_leaf_20_clk),
    .D(net427),
    .RESET_B(net293),
    .SCD(clknet_1_1__leaf_net449),
    .SCE(net446),
    .SET_B(net296),
    .Q(net457),
    .Q_N(net456));
 sky130_fd_sc_hd__sdfxbp_1 c451 (.CLK(clknet_leaf_20_clk),
    .D(net934),
    .SCD(clknet_1_1__leaf_net449),
    .SCE(net863),
    .Q(net459),
    .Q_N(net458));
 sky130_fd_sc_hd__sdfxbp_1 c452 (.CLK(clknet_leaf_20_clk),
    .D(net315),
    .SCD(net455),
    .SCE(net249),
    .Q(net461),
    .Q_N(net460));
 sky130_fd_sc_hd__and3_1 c453 (.A(net461),
    .B(net197),
    .C(net326),
    .X(net462));
 sky130_fd_sc_hd__a2111o_1 c454 (.A1(clknet_1_0__leaf_net432),
    .A2(net440),
    .B1(clknet_1_0__leaf_net287),
    .C1(net293),
    .D1(net458),
    .X(net463));
 sky130_fd_sc_hd__a2111o_1 c455 (.A1(net323),
    .A2(net462),
    .B1(net164),
    .C1(net460),
    .D1(net326),
    .X(net464));
 sky130_fd_sc_hd__sdfbbp_1 c456 (.CLK(clknet_leaf_20_clk),
    .D(net310),
    .RESET_B(net456),
    .SCD(clknet_1_1__leaf_net463),
    .SCE(net985),
    .SET_B(clknet_1_0__leaf_net449),
    .Q(net466),
    .Q_N(net465));
 sky130_fd_sc_hd__sdfbbn_1 c457 (.CLK_N(clknet_leaf_20_clk),
    .D(net447),
    .RESET_B(net461),
    .SCD(net450),
    .SCE(clknet_1_0__leaf_net463),
    .SET_B(net465),
    .Q(net467));
 sky130_fd_sc_hd__sdfxtp_2 c458 (.CLK(clknet_leaf_20_clk),
    .D(clknet_1_0__leaf_net463),
    .SCD(net464),
    .SCE(net324),
    .Q(net815));
 sky130_fd_sc_hd__sdfbbn_1 c459 (.CLK_N(clknet_leaf_20_clk),
    .D(net911),
    .RESET_B(net892),
    .SCD(net461),
    .SCE(clknet_1_1__leaf_net463),
    .SET_B(net453),
    .Q(net468));
 sky130_fd_sc_hd__and2_1 c46 (.A(net796),
    .B(net17),
    .X(net21));
 sky130_fd_sc_hd__sdfxtp_1 c460 (.CLK(clknet_leaf_20_clk),
    .D(clknet_1_0__leaf_net449),
    .SCD(net466),
    .SCE(clknet_1_1__leaf_net463),
    .Q(net469));
 sky130_fd_sc_hd__a2111o_1 c461 (.A1(net469),
    .A2(net284),
    .B1(net815),
    .C1(net460),
    .D1(net385),
    .X(net817));
 sky130_fd_sc_hd__or4bb_1 c462 (.A(net206),
    .B(net836),
    .C_N(net815),
    .D_N(net67),
    .X(net470));
 sky130_fd_sc_hd__and3_4 c463 (.A(net211),
    .B(net830),
    .C(net820),
    .X(net822));
 sky130_fd_sc_hd__sdfbbp_1 c464 (.CLK(clknet_leaf_22_clk),
    .D(net375),
    .RESET_B(net983),
    .SCD(net451),
    .SCE(net833),
    .SET_B(net331),
    .Q(net472),
    .Q_N(net471));
 sky130_fd_sc_hd__a2111o_1 c465 (.A1(net329),
    .A2(net438),
    .B1(net138),
    .C1(net5),
    .D1(net940),
    .X(net473));
 sky130_fd_sc_hd__or4bb_1 c466 (.A(net381),
    .B(net836),
    .C_N(net789),
    .D_N(net210),
    .X(net474));
 sky130_fd_sc_hd__sdfxtp_1 c467 (.CLK(clknet_leaf_22_clk),
    .D(net76),
    .SCD(net344),
    .SCE(net77),
    .Q(net475));
 sky130_fd_sc_hd__dfsbp_1 c468 (.CLK(clknet_leaf_18_clk),
    .D(net474),
    .SET_B(net928),
    .Q(net825));
 sky130_fd_sc_hd__and2_0 c469 (.A(net970),
    .B(net145),
    .X(net476));
 sky130_fd_sc_hd__clkbuf_2 c47 (.A(net17),
    .X(net22));
 sky130_fd_sc_hd__dfbbn_1 c470 (.CLK_N(clknet_leaf_18_clk),
    .D(net476),
    .RESET_B(net439),
    .SET_B(net474),
    .Q(net478),
    .Q_N(net477));
 sky130_fd_sc_hd__and2_0 c471 (.A(net335),
    .B(net834),
    .X(net479));
 sky130_fd_sc_hd__and2_1 c472 (.A(net963),
    .B(net840),
    .X(net480));
 sky130_fd_sc_hd__dfsbp_1 c473 (.CLK(clknet_leaf_18_clk),
    .D(net900),
    .SET_B(net480),
    .Q(net481));
 sky130_fd_sc_hd__sdfbbn_1 c474 (.CLK_N(clknet_leaf_22_clk),
    .D(net331),
    .RESET_B(net77),
    .SCD(net822),
    .SCE(net351),
    .SET_B(net910),
    .Q(net483),
    .Q_N(net482));
 sky130_fd_sc_hd__dfbbn_1 c475 (.CLK_N(clknet_leaf_18_clk),
    .D(net925),
    .RESET_B(net470),
    .SET_B(net296),
    .Q(net484));
 sky130_fd_sc_hd__and3_1 c476 (.A(net996),
    .B(net481),
    .C(net478),
    .X(net485));
 sky130_fd_sc_hd__dfstp_1 c477 (.CLK(clknet_leaf_18_clk),
    .D(net473),
    .SET_B(net478),
    .Q(net486));
 sky130_fd_sc_hd__dfbbp_1 c478 (.CLK(clknet_leaf_22_clk),
    .D(net479),
    .RESET_B(net340),
    .SET_B(net839),
    .Q(net487));
 sky130_fd_sc_hd__or4bb_1 c479 (.A(net487),
    .B(net484),
    .C_N(net485),
    .D_N(net477),
    .X(net488));
 sky130_fd_sc_hd__and2_0 c48 (.A(net20),
    .B(net13),
    .X(net23));
 sky130_fd_sc_hd__sdfxbp_1 c480 (.CLK(clknet_leaf_17_clk),
    .D(net485),
    .SCD(net833),
    .SCE(net381),
    .Q(net490),
    .Q_N(net489));
 sky130_fd_sc_hd__sdfxbp_1 c481 (.CLK(clknet_leaf_18_clk),
    .D(net480),
    .SCD(net930),
    .SCE(net822),
    .Q(net492),
    .Q_N(net491));
 sky130_fd_sc_hd__or4bb_1 c482 (.A(net488),
    .B(net492),
    .C_N(net477),
    .D_N(net489),
    .X(net493));
 sky130_fd_sc_hd__and3_1 c487 (.A(clknet_1_0__leaf_net356),
    .B(net824),
    .C(net102),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_1 c488 (.A(net749),
    .X(net495));
 sky130_fd_sc_hd__and3_1 c489 (.A(net240),
    .B(net205),
    .C(net817),
    .X(net496));
 sky130_fd_sc_hd__and2_1 c49 (.A(net18),
    .B(net19),
    .X(net24));
 sky130_fd_sc_hd__and2_1 c490 (.A(net205),
    .B(net811),
    .X(net827));
 sky130_fd_sc_hd__and3_1 c491 (.A(net224),
    .B(net138),
    .C(net815),
    .X(net497));
 sky130_fd_sc_hd__sdfrtp_1 c492 (.CLK(clknet_leaf_24_clk),
    .D(net366),
    .RESET_B(net850),
    .SCD(net216),
    .SCE(net809),
    .Q(net498));
 sky130_fd_sc_hd__sdfxtp_1 c493 (.CLK(clknet_leaf_22_clk),
    .D(net497),
    .SCD(net496),
    .SCE(net944),
    .Q(net499));
 sky130_fd_sc_hd__and3_1 c494 (.A(net472),
    .B(net55),
    .C(net766),
    .X(net500));
 sky130_fd_sc_hd__sdfxtp_1 c495 (.CLK(clknet_leaf_21_clk),
    .D(net327),
    .SCD(net811),
    .SCE(net830),
    .Q(net501));
 sky130_fd_sc_hd__and3_1 c496 (.A(net372),
    .B(net491),
    .C(net811),
    .X(net502));
 sky130_fd_sc_hd__sdfxtp_1 c497 (.CLK(clknet_leaf_25_clk),
    .D(net495),
    .SCD(net494),
    .SCE(net924),
    .Q(net503));
 sky130_fd_sc_hd__and2_0 c498 (.A(net230),
    .B(net498),
    .X(net504));
 sky130_fd_sc_hd__clkbuf_1 c499 (.A(net946),
    .X(net505));
 sky130_fd_sc_hd__buf_2 c50 (.A(in10),
    .X(net25));
 sky130_fd_sc_hd__and3_1 c500 (.A(net503),
    .B(clknet_1_0__leaf_net242),
    .C(net822),
    .X(net506));
 sky130_fd_sc_hd__dfbbn_1 c501 (.CLK_N(clknet_leaf_23_clk),
    .D(net501),
    .RESET_B(net362),
    .SET_B(net505),
    .Q(net507));
 sky130_fd_sc_hd__dfbbn_1 c502 (.CLK_N(clknet_leaf_26_clk),
    .D(net238),
    .RESET_B(net504),
    .SET_B(net506),
    .Q(net832));
 sky130_fd_sc_hd__and3_1 c503 (.A(net500),
    .B(net507),
    .C(net788),
    .X(net823));
 sky130_fd_sc_hd__and2_4 c504 (.A(net108),
    .B(net386),
    .X(net508));
 sky130_fd_sc_hd__dfstp_2 c505 (.CLK(clknet_leaf_3_clk),
    .D(net114),
    .SET_B(net508),
    .Q(net509));
 sky130_fd_sc_hd__dfstp_1 c506 (.CLK(clknet_leaf_5_clk),
    .D(net508),
    .SET_B(net808),
    .Q(net510));
 sky130_fd_sc_hd__dlrbn_1 c507 (.D(net938),
    .GATE_N(clknet_leaf_5_clk),
    .RESET_B(net508),
    .Q(net511));
 sky130_fd_sc_hd__and2_0 c508 (.A(net392),
    .B(net768),
    .X(net512));
 sky130_fd_sc_hd__and2_0 c509 (.A(net511),
    .B(net512),
    .X(net513));
 sky130_fd_sc_hd__buf_2 c51 (.A(net873),
    .X(net26));
 sky130_fd_sc_hd__and2_0 c510 (.A(net107),
    .B(net512),
    .X(net514));
 sky130_fd_sc_hd__dlrbn_1 c511 (.D(net513),
    .GATE_N(clknet_leaf_5_clk),
    .RESET_B(clknet_1_1__leaf_net260),
    .Q(net515));
 sky130_fd_sc_hd__and2_1 c512 (.A(net386),
    .B(net938),
    .X(net516));
 sky130_fd_sc_hd__and3_1 c513 (.A(net393),
    .B(clknet_1_1__leaf_net253),
    .C(net510),
    .X(net517));
 sky130_fd_sc_hd__dlrbp_1 c514 (.D(clknet_1_1__leaf_net255),
    .GATE(clknet_leaf_11_clk),
    .RESET_B(net387),
    .Q(net519),
    .Q_N(net518));
 sky130_fd_sc_hd__and2_0 c515 (.A(net512),
    .B(net768),
    .X(net520));
 sky130_fd_sc_hd__dlrbp_1 c516 (.D(net112),
    .GATE(clknet_leaf_3_clk),
    .RESET_B(net107),
    .Q(net521));
 sky130_fd_sc_hd__dlrtn_1 c517 (.D(clknet_1_0__leaf_net253),
    .GATE_N(clknet_leaf_9_clk),
    .RESET_B(net516),
    .Q(net522));
 sky130_fd_sc_hd__and2_0 c518 (.A(net522),
    .B(net768),
    .X(net523));
 sky130_fd_sc_hd__and3_1 c519 (.A(net521),
    .B(net509),
    .C(net522),
    .X(net524));
 sky130_fd_sc_hd__and2_1 c52 (.A(net24),
    .B(net22),
    .X(net27));
 sky130_fd_sc_hd__dlrtn_1 c520 (.D(clknet_1_0__leaf_net517),
    .GATE_N(clknet_leaf_9_clk),
    .RESET_B(clknet_1_1__leaf_net253),
    .Q(net525));
 sky130_fd_sc_hd__dlrtn_2 c521 (.D(net514),
    .GATE_N(clknet_leaf_7_clk),
    .RESET_B(net522),
    .Q(net526));
 sky130_fd_sc_hd__dlrtp_1 c522 (.D(net520),
    .GATE(clknet_leaf_4_clk),
    .RESET_B(net508),
    .Q(net527));
 sky130_fd_sc_hd__dfbbp_1 c523 (.CLK(clknet_leaf_9_clk),
    .D(net525),
    .RESET_B(net526),
    .SET_B(clknet_1_1__leaf_net517),
    .Q(net529),
    .Q_N(net528));
 sky130_fd_sc_hd__and2_0 c524 (.A(net515),
    .B(net510),
    .X(net530));
 sky130_fd_sc_hd__and2_0 c525 (.A(net804),
    .B(net526),
    .X(net531));
 sky130_fd_sc_hd__and2_0 c526 (.A(net524),
    .B(clknet_1_1__leaf_net252),
    .X(net532));
 sky130_fd_sc_hd__and2_0 c527 (.A(net8),
    .B(net145),
    .X(net533));
 sky130_fd_sc_hd__and2_0 c528 (.A(clknet_1_0__leaf_net252),
    .B(net408),
    .X(net534));
 sky130_fd_sc_hd__and2_0 c529 (.A(net396),
    .B(net800),
    .X(net535));
 sky130_fd_sc_hd__buf_1 c53 (.A(net873),
    .X(net28));
 sky130_fd_sc_hd__and2_0 c530 (.A(net535),
    .B(net378),
    .X(net536));
 sky130_fd_sc_hd__and2_4 c531 (.A(net417),
    .B(net883),
    .X(net537));
 sky130_fd_sc_hd__dlrtp_1 c532 (.D(net117),
    .GATE(clknet_leaf_4_clk),
    .RESET_B(net508),
    .Q(net538));
 sky130_fd_sc_hd__and2_0 c533 (.A(net532),
    .B(net834),
    .X(net539));
 sky130_fd_sc_hd__dlrtp_1 c534 (.D(net394),
    .GATE(clknet_leaf_4_clk),
    .RESET_B(net537),
    .Q(net540));
 sky130_fd_sc_hd__and2_0 c535 (.A(net974),
    .B(net818),
    .X(net541));
 sky130_fd_sc_hd__edfxbp_1 c536 (.CLK(clknet_leaf_10_clk),
    .D(clknet_1_0__leaf_net539),
    .DE(net537),
    .Q(net542));
 sky130_fd_sc_hd__edfxtp_1 c537 (.CLK(clknet_leaf_9_clk),
    .D(net533),
    .DE(net526),
    .Q(net543));
 sky130_fd_sc_hd__sdlclkp_1 c538 (.CLK(clknet_leaf_7_clk),
    .GATE(net891),
    .SCE(net537),
    .GCLK(net544));
 sky130_fd_sc_hd__and2_2 c539 (.A(net415),
    .B(net540),
    .X(net545));
 sky130_fd_sc_hd__dfbbn_1 c54 (.CLK_N(clknet_leaf_35_clk),
    .D(net795),
    .RESET_B(net22),
    .SET_B(net27),
    .Q(net30),
    .Q_N(net29));
 sky130_fd_sc_hd__and2_0 c540 (.A(net523),
    .B(net545),
    .X(net546));
 sky130_fd_sc_hd__sdlclkp_2 c541 (.CLK(clknet_leaf_10_clk),
    .GATE(net541),
    .SCE(clknet_1_1__leaf_net539),
    .GCLK(net547));
 sky130_fd_sc_hd__sdlclkp_4 c542 (.CLK(clknet_leaf_10_clk),
    .GATE(net546),
    .SCE(net537),
    .GCLK(net814));
 sky130_fd_sc_hd__sdfxbp_1 c543 (.CLK(clknet_leaf_7_clk),
    .D(net403),
    .SCD(net546),
    .SCE(clknet_1_1__leaf_net814),
    .Q(net548));
 sky130_fd_sc_hd__mux4_1 c544 (.A0(net547),
    .A1(net548),
    .A2(net533),
    .A3(net403),
    .S0(clknet_1_1__leaf_net252),
    .S1(net537),
    .X(net549));
 sky130_fd_sc_hd__sdfrtp_1 c545 (.CLK(clknet_leaf_10_clk),
    .D(net534),
    .RESET_B(net884),
    .SCD(clknet_1_0__leaf_net814),
    .SCE(net262),
    .Q(net550));
 sky130_fd_sc_hd__and3_1 c546 (.A(net436),
    .B(net26),
    .C(net518),
    .X(net551));
 sky130_fd_sc_hd__sdfxbp_1 c547 (.CLK(clknet_leaf_9_clk),
    .D(net26),
    .SCD(net508),
    .SCE(net937),
    .Q(net553),
    .Q_N(net552));
 sky130_fd_sc_hd__and2_2 c548 (.A(net551),
    .B(net865),
    .X(net554));
 sky130_fd_sc_hd__sdfxtp_1 c549 (.CLK(clknet_leaf_11_clk),
    .D(net267),
    .SCD(net420),
    .SCE(net554),
    .Q(net555));
 sky130_fd_sc_hd__clkbuf_1 c55 (.A(net30),
    .X(net31));
 sky130_fd_sc_hd__sdfbbn_1 c550 (.CLK_N(clknet_leaf_1_clk),
    .D(net531),
    .RESET_B(net962),
    .SCD(clknet_1_0__leaf_net814),
    .SCE(net121),
    .SET_B(net380),
    .Q(net556));
 sky130_fd_sc_hd__and3_1 c551 (.A(net556),
    .B(clknet_1_1__leaf_net165),
    .C(clknet_1_0__leaf_net814),
    .X(net557));
 sky130_fd_sc_hd__and3_1 c552 (.A(net301),
    .B(net5),
    .C(net770),
    .X(net558));
 sky130_fd_sc_hd__and3_1 c553 (.A(net554),
    .B(net138),
    .C(clknet_1_1__leaf_net757),
    .X(net559));
 sky130_fd_sc_hd__and3_1 c554 (.A(net420),
    .B(net440),
    .C(net552),
    .X(net560));
 sky130_fd_sc_hd__clkbuf_1 c555 (.A(net734),
    .X(net561));
 sky130_fd_sc_hd__and2_0 c556 (.A(net791),
    .B(net419),
    .X(net821));
 sky130_fd_sc_hd__and2_1 c557 (.A(net262),
    .B(net436),
    .X(net562));
 sky130_fd_sc_hd__sdfxtp_1 c558 (.CLK(clknet_leaf_11_clk),
    .D(net557),
    .SCD(net791),
    .SCE(net811),
    .Q(net563));
 sky130_fd_sc_hd__and2_2 c559 (.A(net560),
    .B(net526),
    .X(net564));
 sky130_fd_sc_hd__and3_1 c56 (.A(net799),
    .B(net28),
    .C(net25),
    .X(net32));
 sky130_fd_sc_hd__and2_0 c560 (.A(net264),
    .B(net788),
    .X(net565));
 sky130_fd_sc_hd__buf_1 c561 (.A(net734),
    .X(net566));
 sky130_fd_sc_hd__and3_1 c562 (.A(net561),
    .B(net564),
    .C(net988),
    .X(net567));
 sky130_fd_sc_hd__dfrbp_1 c563 (.CLK(clknet_leaf_11_clk),
    .D(net567),
    .RESET_B(net866),
    .Q(net569),
    .Q_N(net568));
 sky130_fd_sc_hd__mux4_1 c564 (.A0(net569),
    .A1(net379),
    .A2(net564),
    .A3(net554),
    .S0(net115),
    .S1(net508),
    .X(net570));
 sky130_fd_sc_hd__and3_1 c565 (.A(net301),
    .B(net563),
    .C(net568),
    .X(net571));
 sky130_fd_sc_hd__and2_4 c566 (.A(net571),
    .B(net569),
    .X(net572));
 sky130_fd_sc_hd__buf_2 c567 (.A(net724),
    .X(net573));
 sky130_fd_sc_hd__a2111o_1 c568 (.A1(net164),
    .A2(net408),
    .B1(net573),
    .C1(net828),
    .D1(net815),
    .X(net574));
 sky130_fd_sc_hd__and2_0 c569 (.A(net542),
    .B(net550),
    .X(net575));
 sky130_fd_sc_hd__and2_1 c57 (.A(net31),
    .B(net29),
    .X(net33));
 sky130_fd_sc_hd__and3_1 c570 (.A(net429),
    .B(net573),
    .C(net770),
    .X(net576));
 sky130_fd_sc_hd__and3_1 c571 (.A(net387),
    .B(net573),
    .C(net576),
    .X(net577));
 sky130_fd_sc_hd__buf_1 c572 (.A(net724),
    .X(net578));
 sky130_fd_sc_hd__a2111o_4 c573 (.A1(net562),
    .A2(net835),
    .B1(net428),
    .C1(net578),
    .D1(net764),
    .X(net579));
 sky130_fd_sc_hd__mux4_1 c574 (.A0(net519),
    .A1(net578),
    .A2(net121),
    .A3(net408),
    .S0(net573),
    .S1(net579),
    .X(net580));
 sky130_fd_sc_hd__and2_0 c575 (.A(net544),
    .B(net575),
    .X(net581));
 sky130_fd_sc_hd__sdfxtp_1 c576 (.CLK(clknet_leaf_19_clk),
    .D(net408),
    .SCD(net926),
    .SCE(net324),
    .Q(net582));
 sky130_fd_sc_hd__mux4_1 c577 (.A0(net450),
    .A1(net830),
    .A2(net578),
    .A3(net579),
    .S0(net573),
    .S1(net769),
    .X(net583));
 sky130_fd_sc_hd__and3_1 c578 (.A(net284),
    .B(net576),
    .C(net815),
    .X(net584));
 sky130_fd_sc_hd__mux4_1 c579 (.A0(net584),
    .A1(net578),
    .A2(net387),
    .A3(net579),
    .S0(net833),
    .S1(net576),
    .X(net585));
 sky130_fd_sc_hd__dfrbp_1 c58 (.CLK(clknet_leaf_35_clk),
    .D(net17),
    .RESET_B(net14),
    .Q(net35),
    .Q_N(net34));
 sky130_fd_sc_hd__and2_0 c580 (.A(net448),
    .B(net776),
    .X(net586));
 sky130_fd_sc_hd__and2_0 c581 (.A(net377),
    .B(net550),
    .X(net587));
 sky130_fd_sc_hd__and3_1 c582 (.A(net454),
    .B(net566),
    .C(net815),
    .X(net588));
 sky130_fd_sc_hd__and2_0 c583 (.A(net543),
    .B(net775),
    .X(net589));
 sky130_fd_sc_hd__and3_1 c584 (.A(net555),
    .B(net586),
    .C(net566),
    .X(net590));
 sky130_fd_sc_hd__dfbbn_1 c585 (.CLK_N(clknet_leaf_13_clk),
    .D(net587),
    .RESET_B(net584),
    .SET_B(net774),
    .Q(net591));
 sky130_fd_sc_hd__and3_1 c586 (.A(net576),
    .B(net591),
    .C(net573),
    .X(net592));
 sky130_fd_sc_hd__and3_1 c587 (.A(net589),
    .B(net576),
    .C(net592),
    .X(net593));
 sky130_fd_sc_hd__dfbbn_1 c588 (.CLK_N(clknet_leaf_13_clk),
    .D(net989),
    .RESET_B(net593),
    .SET_B(net55),
    .Q(net595),
    .Q_N(net594));
 sky130_fd_sc_hd__and3_1 c589 (.A(net490),
    .B(net67),
    .C(clknet_1_1__leaf_net814),
    .X(net596));
 sky130_fd_sc_hd__and3_2 c59 (.A(net33),
    .B(net22),
    .C(net31),
    .X(net36));
 sky130_fd_sc_hd__dfbbp_1 c590 (.CLK(clknet_leaf_18_clk),
    .D(net77),
    .RESET_B(net880),
    .SET_B(net951),
    .Q(net597));
 sky130_fd_sc_hd__sdfxbp_1 c591 (.CLK(clknet_leaf_19_clk),
    .D(net508),
    .SCD(clknet_1_0__leaf_net596),
    .SCE(net828),
    .Q(net598));
 sky130_fd_sc_hd__and3_1 c592 (.A(net429),
    .B(net598),
    .C(net582),
    .X(net599));
 sky130_fd_sc_hd__and3_4 c593 (.A(net175),
    .B(net572),
    .C(net348),
    .X(net600));
 sky130_fd_sc_hd__or4bb_2 c594 (.A(net344),
    .B(net352),
    .C_N(net838),
    .D_N(net829),
    .X(net601));
 sky130_fd_sc_hd__mux4_1 c595 (.A0(net566),
    .A1(net581),
    .A2(net349),
    .A3(net428),
    .S0(net841),
    .S1(net831),
    .X(net602));
 sky130_fd_sc_hd__sdfbbp_1 c596 (.CLK(clknet_leaf_19_clk),
    .D(net330),
    .RESET_B(net378),
    .SCD(net822),
    .SCE(net428),
    .SET_B(net482),
    .Q(net603));
 sky130_fd_sc_hd__sdfxbp_1 c597 (.CLK(clknet_leaf_19_clk),
    .D(net600),
    .SCD(net603),
    .SCE(net837),
    .Q(net605),
    .Q_N(net604));
 sky130_fd_sc_hd__mux4_1 c598 (.A0(net788),
    .A1(net347),
    .A2(net600),
    .A3(net604),
    .S0(net594),
    .S1(net216),
    .X(net606));
 sky130_fd_sc_hd__sdfrtp_1 c599 (.CLK(clknet_leaf_17_clk),
    .D(net349),
    .RESET_B(net882),
    .SCD(net249),
    .SCE(net526),
    .Q(net607));
 sky130_fd_sc_hd__dfbbp_1 c60 (.CLK(clknet_leaf_33_clk),
    .D(net27),
    .RESET_B(net33),
    .SET_B(net28),
    .Q(net38),
    .Q_N(net37));
 sky130_fd_sc_hd__sdfsbp_1 c600 (.CLK(clknet_leaf_17_clk),
    .D(net529),
    .SCD(net446),
    .SCE(net842),
    .SET_B(net885),
    .Q(net819));
 sky130_fd_sc_hd__and3_1 c601 (.A(net582),
    .B(net599),
    .C(net605),
    .X(net608));
 sky130_fd_sc_hd__sdfxtp_1 c602 (.CLK(clknet_leaf_18_clk),
    .D(clknet_1_1__leaf_net287),
    .SCD(net597),
    .SCE(net601),
    .Q(net609));
 sky130_fd_sc_hd__and3_1 c603 (.A(net346),
    .B(net764),
    .C(net778),
    .X(net610));
 sky130_fd_sc_hd__sdfxtp_1 c604 (.CLK(clknet_leaf_19_clk),
    .D(net347),
    .SCD(net590),
    .SCE(net608),
    .Q(net611));
 sky130_fd_sc_hd__sdfsbp_1 c605 (.CLK(clknet_leaf_17_clk),
    .D(net608),
    .SCD(net904),
    .SCE(net935),
    .SET_B(net882),
    .Q(net816));
 sky130_fd_sc_hd__or4bb_1 c606 (.A(net526),
    .B(net610),
    .C_N(net611),
    .D_N(clknet_1_1__leaf_net596),
    .X(net612));
 sky130_fd_sc_hd__sdfbbn_1 c607 (.CLK_N(clknet_leaf_17_clk),
    .D(net929),
    .RESET_B(net600),
    .SCD(net608),
    .SCE(net822),
    .SET_B(net777),
    .Q(net614),
    .Q_N(net613));
 sky130_fd_sc_hd__sdfxtp_1 c608 (.CLK(clknet_leaf_17_clk),
    .D(net896),
    .SCD(net612),
    .SCE(net992),
    .Q(net615));
 sky130_fd_sc_hd__and3_1 c61 (.A(net952),
    .B(net24),
    .C(net33),
    .X(net39));
 sky130_fd_sc_hd__dfrbp_1 c62 (.CLK(clknet_leaf_35_clk),
    .D(net39),
    .RESET_B(net853),
    .Q(net41),
    .Q_N(net40));
 sky130_fd_sc_hd__and2_0 c63 (.A(net41),
    .B(net21),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 c630 (.A(net117),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_1 c631 (.A(net740),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_1 c632 (.A(net740),
    .X(net618));
 sky130_fd_sc_hd__dfrbp_1 c633 (.CLK(clknet_leaf_7_clk),
    .D(net376),
    .RESET_B(net380),
    .Q(net620),
    .Q_N(net619));
 sky130_fd_sc_hd__and2_0 c634 (.A(net120),
    .B(net509),
    .X(net621));
 sky130_fd_sc_hd__buf_1 c635 (.A(net617),
    .X(net622));
 sky130_fd_sc_hd__buf_1 c636 (.A(net785),
    .X(net623));
 sky130_fd_sc_hd__and2_0 c637 (.A(net623),
    .B(net376),
    .X(net624));
 sky130_fd_sc_hd__and2_0 c638 (.A(net262),
    .B(net623),
    .X(net625));
 sky130_fd_sc_hd__and2_0 c639 (.A(net621),
    .B(net623),
    .X(net626));
 sky130_fd_sc_hd__and2_1 c64 (.A(net38),
    .B(net793),
    .X(net43));
 sky130_fd_sc_hd__and2_0 c640 (.A(net626),
    .B(net620),
    .X(net627));
 sky130_fd_sc_hd__and2_0 c641 (.A(net243),
    .B(net617),
    .X(net628));
 sky130_fd_sc_hd__dfrtn_1 c642 (.CLK_N(clknet_leaf_8_clk),
    .D(net627),
    .RESET_B(net623),
    .Q(net629));
 sky130_fd_sc_hd__clkbuf_1 c643 (.A(net625),
    .X(net630));
 sky130_fd_sc_hd__dfrtp_1 c644 (.CLK(clknet_leaf_5_clk),
    .D(net808),
    .RESET_B(net630),
    .Q(net631));
 sky130_fd_sc_hd__dfrtp_1 c645 (.CLK(clknet_leaf_8_clk),
    .D(net627),
    .RESET_B(net854),
    .Q(net632));
 sky130_fd_sc_hd__and3_2 c646 (.A(net616),
    .B(net632),
    .C(net631),
    .X(net633));
 sky130_fd_sc_hd__and2_0 c647 (.A(net631),
    .B(net628),
    .X(net634));
 sky130_fd_sc_hd__dfrtp_1 c648 (.CLK(clknet_leaf_5_clk),
    .D(net630),
    .RESET_B(net848),
    .Q(net635));
 sky130_fd_sc_hd__or4bb_1 c649 (.A(net392),
    .B(net635),
    .C_N(net633),
    .D_N(net632),
    .X(net636));
 sky130_fd_sc_hd__buf_1 c65 (.A(net19),
    .X(net44));
 sky130_fd_sc_hd__a2111o_1 c650 (.A1(net905),
    .A2(net509),
    .B1(net621),
    .C1(net633),
    .D1(net379),
    .X(net637));
 sky130_fd_sc_hd__and2_0 c651 (.A(net807),
    .B(net624),
    .X(net638));
 sky130_fd_sc_hd__dfsbp_1 c652 (.CLK(clknet_leaf_6_clk),
    .D(net530),
    .SET_B(net421),
    .Q(net640),
    .Q_N(net639));
 sky130_fd_sc_hd__dfsbp_1 c653 (.CLK(clknet_leaf_6_clk),
    .D(net638),
    .SET_B(net867),
    .Q(net641));
 sky130_fd_sc_hd__and2_1 c654 (.A(net618),
    .B(net144),
    .X(net642));
 sky130_fd_sc_hd__and2_2 c655 (.A(net641),
    .B(net906),
    .X(net643));
 sky130_fd_sc_hd__and2_1 c656 (.A(net624),
    .B(net633),
    .X(net644));
 sky130_fd_sc_hd__sdfbbn_1 c657 (.CLK_N(clknet_leaf_6_clk),
    .D(net536),
    .RESET_B(net642),
    .SCD(net636),
    .SCE(net379),
    .SET_B(net545),
    .Q(net645));
 sky130_fd_sc_hd__dfstp_1 c658 (.CLK(clknet_leaf_7_clk),
    .D(net276),
    .SET_B(net643),
    .Q(net646));
 sky130_fd_sc_hd__dfstp_1 c659 (.CLK(clknet_leaf_8_clk),
    .D(net644),
    .SET_B(net869),
    .Q(net647));
 sky130_fd_sc_hd__and2_1 c66 (.A(net2),
    .B(net10),
    .X(net45));
 sky130_fd_sc_hd__and2_1 c660 (.A(net975),
    .B(net631),
    .X(net648));
 sky130_fd_sc_hd__dfstp_1 c661 (.CLK(clknet_leaf_7_clk),
    .D(net421),
    .SET_B(net637),
    .Q(net649));
 sky130_fd_sc_hd__and2_0 c662 (.A(net538),
    .B(net648),
    .X(net650));
 sky130_fd_sc_hd__sdfstp_1 c663 (.CLK(clknet_leaf_6_clk),
    .D(net634),
    .SCD(net262),
    .SCE(net537),
    .SET_B(net941),
    .Q(net651));
 sky130_fd_sc_hd__sdfbbp_1 c664 (.CLK(clknet_leaf_5_clk),
    .D(net855),
    .RESET_B(net648),
    .SCD(net634),
    .SCE(net115),
    .SET_B(net859),
    .Q(net653),
    .Q_N(net652));
 sky130_fd_sc_hd__and3_1 c665 (.A(net269),
    .B(net650),
    .C(net509),
    .X(net654));
 sky130_fd_sc_hd__dlrbn_1 c666 (.D(net997),
    .GATE_N(clknet_leaf_6_clk),
    .RESET_B(net644),
    .Q(net655));
 sky130_fd_sc_hd__and3_4 c667 (.A(net628),
    .B(net649),
    .C(net652),
    .X(net656));
 sky130_fd_sc_hd__sdfstp_1 c668 (.CLK(clknet_leaf_6_clk),
    .D(net655),
    .SCD(net633),
    .SCE(net656),
    .SET_B(net855),
    .Q(net657));
 sky130_fd_sc_hd__sdfbbn_1 c669 (.CLK_N(clknet_leaf_8_clk),
    .D(net1),
    .RESET_B(net644),
    .SCD(net657),
    .SCE(net656),
    .SET_B(net633),
    .Q(net658));
 sky130_fd_sc_hd__clkbuf_1 c67 (.A(net786),
    .X(net46));
 sky130_fd_sc_hd__dlrbn_1 c670 (.D(net636),
    .GATE_N(clknet_leaf_8_clk),
    .RESET_B(net658),
    .Q(net659));
 sky130_fd_sc_hd__and2_1 c671 (.A(net645),
    .B(net657),
    .X(net660));
 sky130_fd_sc_hd__and2_0 c672 (.A(net554),
    .B(net633),
    .X(net661));
 sky130_fd_sc_hd__dlrbp_1 c673 (.D(net424),
    .GATE(clknet_leaf_9_clk),
    .RESET_B(net537),
    .Q(net662));
 sky130_fd_sc_hd__and3_1 c674 (.A(net545),
    .B(net553),
    .C(net629),
    .X(net663));
 sky130_fd_sc_hd__dlrbp_1 c675 (.D(net889),
    .GATE(clknet_leaf_8_clk),
    .RESET_B(net661),
    .Q(net665),
    .Q_N(net664));
 sky130_fd_sc_hd__and2_0 c676 (.A(net144),
    .B(net545),
    .X(net666));
 sky130_fd_sc_hd__or4bb_1 c677 (.A(net622),
    .B(net665),
    .C_N(net552),
    .D_N(net666),
    .X(net667));
 sky130_fd_sc_hd__mux4_1 c678 (.A0(net663),
    .A1(net26),
    .A2(net667),
    .A3(net440),
    .S0(net380),
    .S1(net564),
    .X(net668));
 sky130_fd_sc_hd__or4bb_2 c679 (.A(net26),
    .B(net642),
    .C_N(net545),
    .D_N(net5),
    .X(net669));
 sky130_fd_sc_hd__clkbuf_1 c68 (.A(net46),
    .X(net47));
 sky130_fd_sc_hd__and3_1 c680 (.A(net984),
    .B(net789),
    .C(net779),
    .X(net670));
 sky130_fd_sc_hd__and3_1 c681 (.A(net646),
    .B(net662),
    .C(net622),
    .X(net671));
 sky130_fd_sc_hd__and3_1 c682 (.A(net653),
    .B(net659),
    .C(net564),
    .X(net672));
 sky130_fd_sc_hd__and3_1 c683 (.A(net379),
    .B(net666),
    .C(net622),
    .X(net673));
 sky130_fd_sc_hd__dfbbn_1 c684 (.CLK_N(clknet_leaf_9_clk),
    .D(clknet_1_1__leaf_net165),
    .RESET_B(net673),
    .SET_B(net669),
    .Q(net674));
 sky130_fd_sc_hd__and3_1 c685 (.A(net5),
    .B(net553),
    .C(net622),
    .X(net675));
 sky130_fd_sc_hd__and2_1 c686 (.A(net648),
    .B(net671),
    .X(net676));
 sky130_fd_sc_hd__dfbbn_1 c687 (.CLK_N(clknet_leaf_9_clk),
    .D(net675),
    .RESET_B(net379),
    .SET_B(net664),
    .Q(net678),
    .Q_N(net677));
 sky130_fd_sc_hd__sdfstp_1 c688 (.CLK(clknet_leaf_8_clk),
    .D(net564),
    .SCD(net554),
    .SCE(net669),
    .SET_B(net780),
    .Q(net679));
 sky130_fd_sc_hd__dlrtn_1 c689 (.D(net654),
    .GATE_N(clknet_leaf_6_clk),
    .RESET_B(net787),
    .Q(net680));
 sky130_fd_sc_hd__dfrtn_1 c69 (.CLK_N(clknet_leaf_34_clk),
    .D(net42),
    .RESET_B(net43),
    .Q(net48));
 sky130_fd_sc_hd__and3_1 c690 (.A(net897),
    .B(net680),
    .C(net26),
    .X(net681));
 sky130_fd_sc_hd__dfbbp_1 c691 (.CLK(clknet_leaf_8_clk),
    .D(net670),
    .RESET_B(net672),
    .SET_B(net681),
    .Q(net683),
    .Q_N(net682));
 sky130_fd_sc_hd__sedfxbp_1 c692 (.CLK(clknet_leaf_9_clk),
    .D(net674),
    .DE(net667),
    .SCD(net948),
    .SCE(net545),
    .Q(net685),
    .Q_N(net684));
 sky130_fd_sc_hd__sdfxbp_1 c693 (.CLK(clknet_leaf_14_clk),
    .D(net637),
    .SCD(net643),
    .SCE(net676),
    .Q(net686));
 sky130_fd_sc_hd__sdfxbp_1 c694 (.CLK(clknet_leaf_14_clk),
    .D(net121),
    .SCD(net683),
    .SCE(net684),
    .Q(net687));
 sky130_fd_sc_hd__sdfxtp_1 c695 (.CLK(clknet_leaf_7_clk),
    .D(net967),
    .SCD(net619),
    .SCE(net121),
    .Q(net688));
 sky130_fd_sc_hd__and3_2 c696 (.A(net685),
    .B(net181),
    .C(net385),
    .X(net689));
 sky130_fd_sc_hd__sdfbbn_1 c697 (.CLK_N(clknet_leaf_14_clk),
    .D(net642),
    .RESET_B(net656),
    .SCD(net689),
    .SCE(net643),
    .SET_B(net509),
    .Q(net690));
 sky130_fd_sc_hd__sdfxtp_1 c698 (.CLK(clknet_leaf_14_clk),
    .D(net558),
    .SCD(net440),
    .SCE(net959),
    .Q(net691));
 sky130_fd_sc_hd__sdfxtp_1 c699 (.CLK(clknet_leaf_14_clk),
    .D(net324),
    .SCD(net678),
    .SCE(net684),
    .Q(net692));
 sky130_fd_sc_hd__clkbuf_2 c70 (.A(net47),
    .X(net49));
 sky130_fd_sc_hd__dlrtn_1 c700 (.D(net689),
    .GATE_N(clknet_leaf_14_clk),
    .RESET_B(net676),
    .Q(net693));
 sky130_fd_sc_hd__and3_1 c701 (.A(net588),
    .B(net691),
    .C(net689),
    .X(net694));
 sky130_fd_sc_hd__and3_1 c702 (.A(net574),
    .B(net592),
    .C(net440),
    .X(net695));
 sky130_fd_sc_hd__dfbbn_1 c703 (.CLK_N(clknet_leaf_14_clk),
    .D(net509),
    .RESET_B(net695),
    .SET_B(net669),
    .Q(net696));
 sky130_fd_sc_hd__dfbbn_1 c704 (.CLK_N(clknet_leaf_14_clk),
    .D(net669),
    .RESET_B(net681),
    .SET_B(net656),
    .Q(net697));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(net380),
    .A1(net690),
    .A2(net677),
    .A3(net660),
    .S0(net689),
    .S1(net643),
    .X(net698));
 sky130_fd_sc_hd__and3_1 c706 (.A(net660),
    .B(net694),
    .C(net138),
    .X(net699));
 sky130_fd_sc_hd__and3_4 c707 (.A(net440),
    .B(net647),
    .C(net683),
    .X(net700));
 sky130_fd_sc_hd__and3_1 c708 (.A(net115),
    .B(net468),
    .C(net700),
    .X(net701));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(net793),
    .A1(net687),
    .A2(net689),
    .A3(net509),
    .S0(net700),
    .S1(net380),
    .X(net702));
 sky130_fd_sc_hd__clkbuf_2 c71 (.A(net728),
    .X(net50));
 sky130_fd_sc_hd__dfbbp_1 c710 (.CLK(clknet_leaf_13_clk),
    .D(net537),
    .RESET_B(net574),
    .SET_B(net857),
    .Q(net703));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net181),
    .A1(net696),
    .A2(net647),
    .A3(net689),
    .S0(net700),
    .S1(net782),
    .X(net704));
 sky130_fd_sc_hd__and3_1 c712 (.A(net800),
    .B(net697),
    .C(net704),
    .X(net705));
 sky130_fd_sc_hd__sdfbbp_1 c713 (.CLK(clknet_leaf_15_clk),
    .D(net705),
    .RESET_B(net887),
    .SCD(net660),
    .SCE(net440),
    .SET_B(net656),
    .Q(net706));
 sky130_fd_sc_hd__a2111o_1 c714 (.A1(net877),
    .A2(net701),
    .B1(net614),
    .C1(net486),
    .D1(net700),
    .X(net707));
 sky130_fd_sc_hd__sedfxbp_1 c715 (.CLK(clknet_leaf_13_clk),
    .D(net249),
    .DE(net452),
    .SCD(net700),
    .SCE(net12),
    .Q(net708));
 sky130_fd_sc_hd__sdfbbn_1 c716 (.CLK_N(clknet_leaf_16_clk),
    .D(net579),
    .RESET_B(net656),
    .SCD(net615),
    .SCE(net700),
    .SET_B(net643),
    .Q(net709));
 sky130_fd_sc_hd__sedfxtp_1 c717 (.CLK(clknet_leaf_13_clk),
    .D(net699),
    .DE(net708),
    .SCD(net579),
    .SCE(net613),
    .Q(net710));
 sky130_fd_sc_hd__sedfxtp_1 c718 (.CLK(clknet_leaf_17_clk),
    .D(net67),
    .DE(net493),
    .SCD(net994),
    .SCE(net579),
    .Q(net711));
 sky130_fd_sc_hd__sdfbbn_1 c719 (.CLK_N(clknet_leaf_16_clk),
    .D(net939),
    .RESET_B(net651),
    .SCD(net8),
    .SCE(net573),
    .SET_B(net579),
    .Q(net712));
 sky130_fd_sc_hd__buf_1 c72 (.A(net32),
    .X(net51));
 sky130_fd_sc_hd__or4bb_1 c720 (.A(net459),
    .B(net710),
    .C_N(net573),
    .D_N(net782),
    .X(net713));
 sky130_fd_sc_hd__sedfxtp_1 c721 (.CLK(clknet_leaf_16_clk),
    .D(net688),
    .DE(net486),
    .SCD(net969),
    .SCE(net579),
    .Q(net714));
 sky130_fd_sc_hd__or4bb_1 c722 (.A(net703),
    .B(net633),
    .C_N(net613),
    .D_N(net773),
    .X(net715));
 sky130_fd_sc_hd__sdfrbp_1 c723 (.CLK(clknet_leaf_15_clk),
    .D(net987),
    .RESET_B(net964),
    .SCD(net614),
    .SCE(net656),
    .Q(net716));
 sky130_fd_sc_hd__sdfrbp_1 c724 (.CLK(clknet_leaf_16_clk),
    .D(net898),
    .RESET_B(net849),
    .SCD(net715),
    .SCE(net781),
    .Q(net717));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net138),
    .A1(net12),
    .A2(net706),
    .A3(net715),
    .S0(net656),
    .S1(net579),
    .X(net718));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net633),
    .A1(net573),
    .A2(net709),
    .A3(net595),
    .S0(net700),
    .S1(net711),
    .X(net719));
 sky130_fd_sc_hd__sdfrtn_1 c727 (.CLK_N(clknet_leaf_15_clk),
    .D(net719),
    .RESET_B(net445),
    .SCD(net643),
    .SCE(net933),
    .Q(net720));
 sky130_fd_sc_hd__or4bb_1 c728 (.A(net711),
    .B(net643),
    .C_N(net720),
    .D_N(net12),
    .X(net721));
 sky130_fd_sc_hd__sdfrtp_1 c729 (.CLK(clknet_leaf_16_clk),
    .D(net721),
    .RESET_B(net878),
    .SCD(net713),
    .SCE(net594),
    .Q(net722));
 sky130_fd_sc_hd__dfrtp_1 c73 (.CLK(clknet_leaf_34_clk),
    .D(net43),
    .RESET_B(net49),
    .Q(net52));
 sky130_fd_sc_hd__and3_1 c730 (.A(net692),
    .B(net722),
    .C(net712),
    .X(net723));
 sky130_fd_sc_hd__or4bb_1 c731 (.A(net693),
    .B(net717),
    .C_N(net723),
    .D_N(net722));
 sky130_fd_sc_hd__buf_1 c74 (.A(net45),
    .X(net53));
 sky130_fd_sc_hd__dfrtp_1 c75 (.CLK(clknet_leaf_34_clk),
    .D(net51),
    .RESET_B(net847),
    .Q(net54));
 sky130_fd_sc_hd__dfrtp_4 c76 (.CLK(clknet_leaf_34_clk),
    .D(net47),
    .RESET_B(net49),
    .Q(net55));
 sky130_fd_sc_hd__sdfrbp_1 c77 (.CLK(clknet_leaf_29_clk),
    .D(net845),
    .RESET_B(net844),
    .SCD(net55),
    .SCE(net53),
    .Q(net57),
    .Q_N(net56));
 sky130_fd_sc_hd__and2_4 c78 (.A(net50),
    .B(net37),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 c79 (.A(net843),
    .X(net59));
 sky130_fd_sc_hd__sdfxbp_1 c80 (.CLK(clknet_leaf_29_clk),
    .D(net48),
    .SCD(net42),
    .SCE(net804),
    .Q(net61),
    .Q_N(net60));
 sky130_fd_sc_hd__and3_1 c81 (.A(net59),
    .B(net58),
    .C(net52),
    .X(net62));
 sky130_fd_sc_hd__and2_1 c82 (.A(net54),
    .B(net40),
    .X(net63));
 sky130_fd_sc_hd__and2_4 c83 (.A(net62),
    .B(net63),
    .X(net831));
 sky130_fd_sc_hd__clkbuf_1 c84 (.A(net981),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 c85 (.A(net915),
    .X(net65));
 sky130_fd_sc_hd__dfsbp_1 c86 (.CLK(clknet_leaf_34_clk),
    .D(net14),
    .SET_B(net18),
    .Q(net66));
 sky130_fd_sc_hd__and2_2 c87 (.A(net789),
    .B(net61),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 c88 (.A(net44),
    .X(net68));
 sky130_fd_sc_hd__dfsbp_1 c89 (.CLK(clknet_leaf_34_clk),
    .D(net893),
    .SET_B(net68),
    .Q(net70),
    .Q_N(net69));
 sky130_fd_sc_hd__dfstp_1 c90 (.CLK(clknet_leaf_34_clk),
    .D(net803),
    .SET_B(net68),
    .Q(net71));
 sky130_fd_sc_hd__and2_1 c91 (.A(net3),
    .B(net5),
    .X(net72));
 sky130_fd_sc_hd__dfstp_1 c92 (.CLK(clknet_leaf_34_clk),
    .D(net18),
    .SET_B(net68),
    .Q(net73));
 sky130_fd_sc_hd__sdfxbp_1 c93 (.CLK(clknet_leaf_27_clk),
    .D(net65),
    .SCD(net67),
    .SCE(net72),
    .Q(net75),
    .Q_N(net74));
 sky130_fd_sc_hd__dfstp_1 c94 (.CLK(clknet_leaf_28_clk),
    .D(net886),
    .SET_B(net68),
    .Q(net76));
 sky130_fd_sc_hd__and2_2 c95 (.A(net76),
    .B(net44),
    .X(net77));
 sky130_fd_sc_hd__and2_0 c96 (.A(net70),
    .B(net75),
    .X(net78));
 sky130_fd_sc_hd__and2_1 c97 (.A(net78),
    .B(net993),
    .X(net79));
 sky130_fd_sc_hd__and3_1 c98 (.A(net63),
    .B(net55),
    .C(net79),
    .X(net80));
 sky130_fd_sc_hd__and2_0 c99 (.A(net73),
    .B(net74),
    .X(net81));
 sky130_fd_sc_hd__sdfrtp_1 merge732 (.CLK(clknet_leaf_13_clk),
    .D(net55),
    .RESET_B(net516),
    .SCD(net577),
    .SCE(net528),
    .Q(net724));
 sky130_fd_sc_hd__sdfrtp_1 merge733 (.CLK(clknet_leaf_32_clk),
    .D(net133),
    .RESET_B(net126),
    .SCE(net135),
    .Q(net154));
 sky130_fd_sc_hd__sdfsbp_1 merge734 (.CLK(clknet_leaf_0_clk),
    .D(net299),
    .SCD(clknet_1_0__leaf_net165),
    .SCE(net413),
    .SET_B(net863),
    .Q(net727),
    .Q_N(net726));
 sky130_fd_sc_hd__dlrtn_1 merge735 (.D(net23),
    .GATE_N(clknet_leaf_34_clk),
    .RESET_B(net53),
    .Q(net728));
 sky130_fd_sc_hd__sdfsbp_1 merge736 (.CLK(clknet_leaf_29_clk),
    .D(net51),
    .SCD(net965),
    .SCE(net788),
    .SET_B(net36),
    .Q(net730),
    .Q_N(net729));
 sky130_fd_sc_hd__sdfbbp_1 merge737 (.CLK(clknet_leaf_36_clk),
    .D(net787),
    .RESET_B(net3),
    .SCD(net9),
    .SCE(net6),
    .SET_B(net11),
    .Q(net732),
    .Q_N(net731));
 sky130_fd_sc_hd__sdfstp_1 merge738 (.CLK(clknet_leaf_2_clk),
    .D(net794),
    .SCD(net111),
    .SCE(net112),
    .SET_B(net808),
    .Q(net733));
 sky130_fd_sc_hd__sdfstp_1 merge739 (.CLK(clknet_leaf_10_clk),
    .D(net559),
    .SCD(net565),
    .SCE(net564),
    .SET_B(net862),
    .Q(net734));
 sky130_fd_sc_hd__sdfxbp_1 merge740 (.CLK(clknet_leaf_28_clk),
    .D(net80),
    .SCD(net93),
    .SCE(net813),
    .Q(net736),
    .Q_N(net735));
 sky130_fd_sc_hd__sdfstp_1 merge741 (.CLK(clknet_leaf_37_clk),
    .D(net917),
    .SCD(net267),
    .SCE(net383),
    .SET_B(net961),
    .Q(net737));
 sky130_fd_sc_hd__sdfxbp_1 merge742 (.CLK(clknet_leaf_4_clk),
    .D(net121),
    .SCD(clknet_1_0__leaf_net255),
    .SCE(clknet_1_0__leaf_net260),
    .Q(net739),
    .Q_N(net738));
 sky130_fd_sc_hd__sdfxtp_1 merge743 (.CLK(clknet_leaf_4_clk),
    .D(clknet_1_1__leaf_net260),
    .SCD(net509),
    .SCE(net382),
    .Q(net740));
 sky130_fd_sc_hd__sdfbbn_1 merge744 (.CLK_N(clknet_leaf_12_clk),
    .D(net309),
    .RESET_B(net121),
    .SCD(net430),
    .SCE(net789),
    .SET_B(net831),
    .Q(net742),
    .Q_N(net741));
 sky130_fd_sc_hd__sdfxtp_1 merge745 (.CLK(clknet_leaf_0_clk),
    .D(clknet_1_1__leaf_net250),
    .SCD(clknet_1_1__leaf_net290),
    .SCE(net147),
    .Q(net743));
 sky130_fd_sc_hd__sedfxbp_1 merge746 (.CLK(clknet_leaf_31_clk),
    .D(net184),
    .DE(net25),
    .SCD(net110),
    .SCE(net249),
    .Q(net745),
    .Q_N(net744));
 sky130_fd_sc_hd__sdfxtp_1 merge747 (.CLK(clknet_leaf_35_clk),
    .D(net24),
    .SCD(net14),
    .SCE(net27),
    .Q(net746));
 sky130_fd_sc_hd__sedfxbp_1 merge748 (.CLK(clknet_leaf_24_clk),
    .D(net214),
    .DE(net82),
    .SCD(net189),
    .SCE(net831),
    .Q(net748),
    .Q_N(net747));
 sky130_fd_sc_hd__sdfbbn_1 merge749 (.CLK_N(clknet_leaf_23_clk),
    .D(net502),
    .RESET_B(net499),
    .SCD(net249),
    .SCE(net829),
    .SET_B(net767),
    .Q(net750),
    .Q_N(net749));
 sky130_fd_sc_hd__dlrtp_1 merge750 (.D(net257),
    .GATE(clknet_leaf_37_clk),
    .RESET_B(net976),
    .Q(net751));
 sky130_fd_sc_hd__dfbbn_1 merge751 (.CLK_N(clknet_leaf_36_clk),
    .D(net9),
    .RESET_B(net127),
    .SET_B(net124),
    .Q(net753),
    .Q_N(net752));
 sky130_fd_sc_hd__dlrtp_1 merge752 (.D(net127),
    .GATE(clknet_leaf_2_clk),
    .RESET_B(clknet_1_0__leaf_net258),
    .Q(net754));
 sky130_fd_sc_hd__dfxtp_1 s753 (.CLK(clknet_leaf_27_clk),
    .D(net84),
    .Q(net755));
 sky130_fd_sc_hd__dfxtp_1 s754 (.CLK(clknet_leaf_37_clk),
    .D(net125),
    .Q(net756));
 sky130_fd_sc_hd__dlclkp_1 s755 (.CLK(clknet_leaf_32_clk),
    .GATE(net168),
    .GCLK(net757));
 sky130_fd_sc_hd__dlclkp_2 s756 (.CLK(clknet_leaf_24_clk),
    .GATE(net241),
    .GCLK(net758));
 sky130_fd_sc_hd__dlclkp_4 s757 (.CLK(clknet_leaf_3_clk),
    .GATE(net263),
    .GCLK(net759));
 sky130_fd_sc_hd__dlxbn_1 s758 (.D(net280),
    .GATE_N(clknet_leaf_38_clk),
    .Q(net761),
    .Q_N(net760));
 sky130_fd_sc_hd__dlxbn_1 s759 (.D(net295),
    .GATE_N(clknet_leaf_0_clk),
    .Q(net762));
 sky130_fd_sc_hd__dlxbp_1 s760 (.D(net307),
    .GATE(clknet_leaf_21_clk),
    .Q(net763));
 sky130_fd_sc_hd__dlxtn_2 s761 (.D(net328),
    .GATE_N(clknet_leaf_20_clk),
    .Q(net764));
 sky130_fd_sc_hd__dlxtn_1 s762 (.D(net370),
    .GATE_N(clknet_leaf_24_clk),
    .Q(net765));
 sky130_fd_sc_hd__dlxtn_1 s763 (.D(net373),
    .GATE_N(clknet_leaf_23_clk),
    .Q(net766));
 sky130_fd_sc_hd__dlxtp_1 s764 (.D(net374),
    .GATE(clknet_leaf_23_clk),
    .Q(net767));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s765 (.D(net388),
    .SLEEP_B(clknet_leaf_10_clk),
    .Q(net768));
 sky130_fd_sc_hd__dfxbp_1 s766 (.CLK(clknet_leaf_12_clk),
    .D(net442),
    .Q(net770),
    .Q_N(net769));
 sky130_fd_sc_hd__dfxbp_1 s767 (.CLK(clknet_leaf_9_clk),
    .D(net549),
    .Q(net772),
    .Q_N(net771));
 sky130_fd_sc_hd__dfxtp_1 s768 (.CLK(clknet_leaf_13_clk),
    .D(net570),
    .Q(net773));
 sky130_fd_sc_hd__dfxtp_1 s769 (.CLK(clknet_leaf_13_clk),
    .D(net580),
    .Q(net774));
 sky130_fd_sc_hd__dfxtp_1 s770 (.CLK(clknet_leaf_13_clk),
    .D(net583),
    .Q(net775));
 sky130_fd_sc_hd__dlclkp_1 s771 (.CLK(clknet_leaf_19_clk),
    .GATE(net585),
    .GCLK(net776));
 sky130_fd_sc_hd__dlclkp_2 s772 (.CLK(clknet_leaf_17_clk),
    .GATE(net602),
    .GCLK(net777));
 sky130_fd_sc_hd__dlclkp_4 s773 (.CLK(clknet_leaf_17_clk),
    .GATE(net606),
    .GCLK(net778));
 sky130_fd_sc_hd__dlxbn_1 s774 (.D(net668),
    .GATE_N(clknet_leaf_8_clk),
    .Q(net780),
    .Q_N(net779));
 sky130_fd_sc_hd__dlxbn_1 s775 (.D(net698),
    .GATE_N(clknet_leaf_15_clk),
    .Q(net782),
    .Q_N(net781));
 sky130_fd_sc_hd__dlxbp_1 s776 (.D(net702),
    .GATE(clknet_leaf_13_clk),
    .Q(net783));
 sky130_fd_sc_hd__dlxtn_1 s777 (.D(net718),
    .GATE_N(clknet_leaf_15_clk),
    .Q(net784));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(in0),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(in1),
    .X(net786));
 sky130_fd_sc_hd__buf_2 input3 (.A(in11),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(in12),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(in13),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(in14),
    .X(net790));
 sky130_fd_sc_hd__buf_2 input7 (.A(in15),
    .X(net791));
 sky130_fd_sc_hd__buf_1 input8 (.A(in16),
    .X(net792));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(in17),
    .X(net793));
 sky130_fd_sc_hd__buf_1 input10 (.A(in18),
    .X(net794));
 sky130_fd_sc_hd__buf_1 input11 (.A(in19),
    .X(net795));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(in2),
    .X(net796));
 sky130_fd_sc_hd__buf_1 input13 (.A(in20),
    .X(net797));
 sky130_fd_sc_hd__buf_1 input14 (.A(in21),
    .X(net798));
 sky130_fd_sc_hd__buf_1 input15 (.A(in22),
    .X(net799));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(in23),
    .X(net800));
 sky130_fd_sc_hd__buf_1 input17 (.A(in24),
    .X(net801));
 sky130_fd_sc_hd__buf_1 input18 (.A(in3),
    .X(net802));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(in4),
    .X(net803));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(in5),
    .X(net804));
 sky130_fd_sc_hd__buf_1 input21 (.A(in6),
    .X(net805));
 sky130_fd_sc_hd__buf_1 input22 (.A(in7),
    .X(net806));
 sky130_fd_sc_hd__buf_1 input23 (.A(in8),
    .X(net807));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(in9),
    .X(net808));
 sky130_fd_sc_hd__buf_2 output25 (.A(net809),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output26 (.A(net810),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output27 (.A(net811),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output28 (.A(net812),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output29 (.A(net813),
    .X(out12));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(clknet_1_1__leaf_net814),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output31 (.A(net815),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output32 (.A(net816),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output33 (.A(net817),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output34 (.A(net818),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output35 (.A(net819),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output36 (.A(net820),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output37 (.A(net821),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output38 (.A(net822),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output39 (.A(net823),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output40 (.A(net824),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output41 (.A(net825),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output42 (.A(net826),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output43 (.A(net827),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output44 (.A(net828),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output45 (.A(net834),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output46 (.A(net830),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output47 (.A(net831),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output48 (.A(net832),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output49 (.A(net833),
    .X(out9));
 sky130_fd_sc_hd__buf_4 fanout50 (.A(net885),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_36_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_37_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_38_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_39_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net390 (.A(net390),
    .X(clknet_0_net390));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net390 (.A(clknet_0_net390),
    .X(clknet_1_0__leaf_net390));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net390 (.A(clknet_0_net390),
    .X(clknet_1_1__leaf_net390));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net757 (.A(net757),
    .X(clknet_0_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net757 (.A(clknet_0_net757),
    .X(clknet_1_0__leaf_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net757 (.A(clknet_0_net757),
    .X(clknet_1_1__leaf_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net814 (.A(net814),
    .X(clknet_0_net814));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net814 (.A(clknet_0_net814),
    .X(clknet_1_0__leaf_net814));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net814 (.A(clknet_0_net814),
    .X(clknet_1_1__leaf_net814));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net596 (.A(net596),
    .X(clknet_0_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net596 (.A(clknet_0_net596),
    .X(clknet_1_0__leaf_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net596 (.A(clknet_0_net596),
    .X(clknet_1_1__leaf_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net432 (.A(net432),
    .X(clknet_0_net432));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net432 (.A(clknet_0_net432),
    .X(clknet_1_0__leaf_net432));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net432 (.A(clknet_0_net432),
    .X(clknet_1_1__leaf_net432));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net463 (.A(net463),
    .X(clknet_0_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net463 (.A(clknet_0_net463),
    .X(clknet_1_0__leaf_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net463 (.A(clknet_0_net463),
    .X(clknet_1_1__leaf_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net261 (.A(net261),
    .X(clknet_0_net261));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net261 (.A(clknet_0_net261),
    .X(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net261 (.A(clknet_0_net261),
    .X(clknet_1_1__leaf_net261));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net399 (.A(net399),
    .X(clknet_0_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_0__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_1__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net402 (.A(net402),
    .X(clknet_0_net402));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net402 (.A(clknet_0_net402),
    .X(clknet_1_0__leaf_net402));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net402 (.A(clknet_0_net402),
    .X(clknet_1_1__leaf_net402));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net398 (.A(net398),
    .X(clknet_0_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_0__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_1__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net401 (.A(net401),
    .X(clknet_0_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net401 (.A(clknet_0_net401),
    .X(clknet_1_0__leaf_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net401 (.A(clknet_0_net401),
    .X(clknet_1_1__leaf_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net250 (.A(net250),
    .X(clknet_0_net250));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net250 (.A(clknet_0_net250),
    .X(clknet_1_0__leaf_net250));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net250 (.A(clknet_0_net250),
    .X(clknet_1_1__leaf_net250));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net287 (.A(net287),
    .X(clknet_0_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net287 (.A(clknet_0_net287),
    .X(clknet_1_0__leaf_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net287 (.A(clknet_0_net287),
    .X(clknet_1_1__leaf_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net449 (.A(net449),
    .X(clknet_0_net449));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net449 (.A(clknet_0_net449),
    .X(clknet_1_0__leaf_net449));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net449 (.A(clknet_0_net449),
    .X(clknet_1_1__leaf_net449));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net258 (.A(net258),
    .X(clknet_0_net258));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net258 (.A(clknet_0_net258),
    .X(clknet_1_0__leaf_net258));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net258 (.A(clknet_0_net258),
    .X(clknet_1_1__leaf_net258));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net252 (.A(net252),
    .X(clknet_0_net252));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net252 (.A(clknet_0_net252),
    .X(clknet_1_0__leaf_net252));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net252 (.A(clknet_0_net252),
    .X(clknet_1_1__leaf_net252));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net539 (.A(net539),
    .X(clknet_0_net539));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net539 (.A(clknet_0_net539),
    .X(clknet_1_0__leaf_net539));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net539 (.A(clknet_0_net539),
    .X(clknet_1_1__leaf_net539));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net253 (.A(net253),
    .X(clknet_0_net253));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net253 (.A(clknet_0_net253),
    .X(clknet_1_0__leaf_net253));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net253 (.A(clknet_0_net253),
    .X(clknet_1_1__leaf_net253));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net517 (.A(net517),
    .X(clknet_0_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net517 (.A(clknet_0_net517),
    .X(clknet_1_0__leaf_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net517 (.A(clknet_0_net517),
    .X(clknet_1_1__leaf_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net255 (.A(net255),
    .X(clknet_0_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net255 (.A(clknet_0_net255),
    .X(clknet_1_0__leaf_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net255 (.A(clknet_0_net255),
    .X(clknet_1_1__leaf_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net251 (.A(net251),
    .X(clknet_0_net251));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net251 (.A(clknet_0_net251),
    .X(clknet_1_0__leaf_net251));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net251 (.A(clknet_0_net251),
    .X(clknet_1_1__leaf_net251));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net290 (.A(net290),
    .X(clknet_0_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net290 (.A(clknet_0_net290),
    .X(clknet_1_0__leaf_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net290 (.A(clknet_0_net290),
    .X(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net260 (.A(net260),
    .X(clknet_0_net260));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net260 (.A(clknet_0_net260),
    .X(clknet_1_0__leaf_net260));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net260 (.A(clknet_0_net260),
    .X(clknet_1_1__leaf_net260));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net242 (.A(net242),
    .X(clknet_0_net242));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net242 (.A(clknet_0_net242),
    .X(clknet_1_0__leaf_net242));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net242 (.A(clknet_0_net242),
    .X(clknet_1_1__leaf_net242));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net356 (.A(net356),
    .X(clknet_0_net356));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net356 (.A(clknet_0_net356),
    .X(clknet_1_0__leaf_net356));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net356 (.A(clknet_0_net356),
    .X(clknet_1_1__leaf_net356));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net359 (.A(net359),
    .X(clknet_0_net359));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net359 (.A(clknet_0_net359),
    .X(clknet_1_0__leaf_net359));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net359 (.A(clknet_0_net359),
    .X(clknet_1_1__leaf_net359));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net160 (.A(net160),
    .X(clknet_0_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net160 (.A(clknet_0_net160),
    .X(clknet_1_0__leaf_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net160 (.A(clknet_0_net160),
    .X(clknet_1_1__leaf_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net165 (.A(net165),
    .X(clknet_0_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net165 (.A(clknet_0_net165),
    .X(clknet_1_0__leaf_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net165 (.A(clknet_0_net165),
    .X(clknet_1_1__leaf_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net294 (.A(net294),
    .X(clknet_0_net294));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net294 (.A(clknet_0_net294),
    .X(clknet_1_0__leaf_net294));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net294 (.A(clknet_0_net294),
    .X(clknet_1_1__leaf_net294));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net166 (.A(net166),
    .X(clknet_0_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net166 (.A(clknet_0_net166),
    .X(clknet_1_0__leaf_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net166 (.A(clknet_0_net166),
    .X(clknet_1_1__leaf_net166));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net158 (.A(net158),
    .X(clknet_0_net158));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net158 (.A(clknet_0_net158),
    .X(clknet_1_0__leaf_net158));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net158 (.A(clknet_0_net158),
    .X(clknet_1_1__leaf_net158));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net171 (.A(net171),
    .X(clknet_0_net171));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net171 (.A(clknet_0_net171),
    .X(clknet_1_0__leaf_net171));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net171 (.A(clknet_0_net171),
    .X(clknet_1_1__leaf_net171));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net175),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net175),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net836),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net836),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net838),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net836),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net600),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net600),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net728),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net50),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net52),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net247),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net41),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net631),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net714),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net240),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net187),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net189),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net34),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net619),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net527),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net755),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net783),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net195),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net538),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net83),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net201),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net771),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net422),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net56),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net769),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net554),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net618),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net100),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net268),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net175),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net179),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net746),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net793),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net321),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net58),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net385),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net707),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net215),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net475),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net337),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net601),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net394),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net537),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net829),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net71),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net686),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net154),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net629),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net193),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net540),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net457),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net54),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net170),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net185),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net609),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net679),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net716),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net748),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net296),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net416),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net202),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net88),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net607),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net632),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net639),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net281),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net157),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net150),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net764),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net467),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net301),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net86),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net118),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net729),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net203),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net283),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net358),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net178),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net149),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net282),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net754),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net281),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(net499),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net478),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net180),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(net196),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net115),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(net483),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(net490),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(net768),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(net355),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(net784),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(net293),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(net605),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(net408),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(net772),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(net510),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(net595),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(net439),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(net509),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(net48),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(net191),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(net471),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(net305),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(net750),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(net199),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(net682),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(net73),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(net383),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(net486),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(net35),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(net342),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(net292),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(net190),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(net132),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(net820),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(net143),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(net685),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(net136),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(net274),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(net419),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(net393),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(net700),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(net60),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(net75),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(net640),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(net228),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(net711),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(net444),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(net220),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(net357),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(net234),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(net405),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(net635),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(net265),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(net57),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(net98),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(net163),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(net308),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(net730),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(net273),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(net55),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(net553),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(net460),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(net338),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(net620),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(net543),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(net146),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(net284),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(net218),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(net393),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(net69),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(net651),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(net74),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(net439),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(net650),
    .X(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c50_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_D (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c35_B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_X (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_B (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_B (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_X (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_SCD (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_D (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_D (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_X (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_RESET_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_X (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_X (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge746_SCD (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_X (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge738_SCD (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_GATE (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_RESET_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_S0 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_D (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_RESET_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_X (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A0 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_D (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_X (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold94_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_SCE (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_S0 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_S1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_X (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_D_N (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_SCE (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_RESET_B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_X (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_C (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_Q (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge744_RESET_B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge742_D (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_SCE (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_D (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_SCE (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_S1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A3 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_X (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_GATE (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_B (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_B (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge733_RESET_B (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_RESET_B (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_SCD (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_GATE (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_SCE (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_D (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_X (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c48_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c39_X (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_RESET_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge733_SCE (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_SET_B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_D (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_SET_B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_X (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_C (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_X (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_D (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_X (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_Q (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A3 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_Q_N (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold155_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_B (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_Q (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge745_SCE (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S0 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_RESET_B (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_D (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_X (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_D (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_RESET_B (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_DE (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_X (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_GCLK (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_Q (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_S1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_SCE (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_X (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold37_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_X (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold18_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge748_SCD (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_RESET_B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_D_N (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_C1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_X (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c48_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c45_X (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_D (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_S0 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_SCD (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_SET_B (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_Q_N (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c54_RESET_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c52_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c47_X (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_C1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold12_A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_X (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge749_SCD (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge746_SCE (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_D (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_SCD (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_SCE (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_SET_B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_SCE (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_RESET_B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_X (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge746_DE (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c56_C (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c50_X (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_D (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_SCE (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_C (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_D (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_B (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c51_X (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_B (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_SCD (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c638_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_SCE (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_SCE (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_S0 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_X (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge741_SCD (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_D (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_D (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_SCD (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_X (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_RESET_B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_D (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_S0 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_D (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_X (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold127_A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_D (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_SCE (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_SCE (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_X (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold89_A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold73_A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_Q (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold156_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_X (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_SET_B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A3 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_X (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net287_A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_X (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_D (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_X (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold100_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_C1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_RESET_B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_SET_B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_Q (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold66_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_SET_B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_SET_B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_Q (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_S0 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_SET_B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_X (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_D (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_SCE (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_SCE (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_RESET_B (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_SET_B (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_SCD (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_X (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A0 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_SCE (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_SET_B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_SET_B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_X (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge736_SET_B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_X (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_D (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_S0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_SCE (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_SCD (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_D (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_B (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_SCE (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_X (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_B (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_D (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_D (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_X (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_X (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_RESET_B (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_B (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_X (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_RESET_B (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c657_SCE (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c650_D1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_B (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_B (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_X (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A0 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_S0 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_RESET_B (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_SET_B (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_SET_B (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_S0 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_X (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_SCE (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_SCD (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_B (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_RESET_B (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_X (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold43_A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_C (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_D1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_SCD (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_Q (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold158_A (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold129_A (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_A (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_C (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_Q (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c32_B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c30_X (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_RESET_B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A3 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_D (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_SCE (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_SCE (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_DE (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_X (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold102_A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_D (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A3 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A2 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_B (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_C (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_B1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_B (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_Q (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_RESET_B (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_D (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_D1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_SCD (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_C (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_X (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold128_A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_B (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_Q_N (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_SCE (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_C (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_SCD (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A3 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_B (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A2 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S0 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A3 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_Q (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_SCD (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_Q_N (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold117_A (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_DE (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_C1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_Q (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_RESET_B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_RESET_B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_X (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_D (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_SCD (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_D_N (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_C1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c31_X (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_D (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_S1 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_SCD (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_RESET_B (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_RESET_B (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_RESET_B (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_D (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_SET_B (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_X (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold107_A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge743_SCD (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A3 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_D (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_SET_B (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_C (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c650_A2 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_B (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_B (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_Q (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold104_A (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_B (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_C (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_Q (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_SCE (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_B (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_DE (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_B (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_RESET_B (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_Q (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold50_A (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_D (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_RESET_B (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_SCE (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S1 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_SCE (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_SCE (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_DE (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_RESET_B (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_X (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_SCE (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_C_N (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_B (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c657_SET_B (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_B (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_X (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold149_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge732_D (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_SCD (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_Q (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_SET_B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold32_A (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_SCD (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A3 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_SCE (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_X (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge739_SCE (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_D (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_C (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_S1 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_B (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_X (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_C_N (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_SCE (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_C (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_B (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_B (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_B1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_X (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_SCE (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_SET_B (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_SCE (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_SCD (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_D (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A3 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A3 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_X (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge737_SCE (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c32_X (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_SCE (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_D (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_SET_B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_B (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_B (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_SET_B (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_SCD (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_B (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c650_C1 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c649_C_N (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_X (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_D (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_SET_B (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c650_X (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_B (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_SCD (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_SET_B (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_S1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_SCE (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_SCD (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c658_SET_B (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_X (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold160_A (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_RESET_B (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_Q (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S0 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_SCE (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_RESET_B (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_SET_B (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_SET_B (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_RESET_B (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_SCE (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_SCE (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_X (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_SCD (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A3 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_X (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_SCD (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_X (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_D (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_B (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_D_N (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_B (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_B (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_D (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_Q (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold130_A (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_SCE (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_SCD (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_D1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S0 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S0 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_C (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_X (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_SCE (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_X (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_D (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_s754_Q (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_B (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_B (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_B (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_Q (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_D (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold76_A (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_s761_Q (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_B (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_D1 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_B (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_D (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_RESET_B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_SCE (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_D (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_SCD (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_RESET_B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c35_C (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_X (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_D_N (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge748_DE (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_D (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_SCE (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A3 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_X (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_D_N (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_X (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_C (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_D (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_B (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge737_D (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_RESET_B (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_SCE (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge736_SCE (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A0 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_B (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_C (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A3 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge744_SCE (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_B (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_C_N (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_B (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_D (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c33_A (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_SCE (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_SCD (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_B1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A2 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold40_A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A0 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_B (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_B (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_D (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_SCD (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_D (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_C (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_C (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_B (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_SCE (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c28_B (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_B (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge738_SET_B (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_D (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_SET_B (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_B (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_output27_A (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_SCE (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_C (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_SCD (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_B (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_X (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_output31_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_C (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_C (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_D1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_C (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_C_N (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_B1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_Q (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_output33_A (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_C (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_X (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_output34_A (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c30_A (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_X (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold123_A (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_output36_A (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_C (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_B (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_Q (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_output38_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_SCE (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_SCD (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_C (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_SCE (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_SCD (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_X (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_output44_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_SCE (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_C1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_B (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_B (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_X (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold51_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge749_SCE (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_D_N (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_X (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_output46_A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_SCE (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_B (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A3 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_C (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_X (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_output47_A (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge748_SCE (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge744_SET_B (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_X (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_RESET_B (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_SCE (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_DE (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_output49_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_SCD (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_SCE (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_D (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_X (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_X (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_B (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_RESET_B (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_B (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_SCD (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_A (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_B (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_SET_B (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_S1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_SCE (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_X (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_X (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_X (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_X (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_SCD (.DIODE(clknet_1_0__leaf_net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_SCD (.DIODE(clknet_1_0__leaf_net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_C (.DIODE(clknet_1_0__leaf_net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net814_X (.DIODE(clknet_1_0__leaf_net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_SCE (.DIODE(clknet_1_1__leaf_net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_C (.DIODE(clknet_1_1__leaf_net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_output30_A (.DIODE(clknet_1_1__leaf_net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net814_X (.DIODE(clknet_1_1__leaf_net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold12_X (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_SCD (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold43_X (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_SET_B (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold51_X (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_SCE (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_D (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold73_X (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold89_X (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_SET_B (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold94_X (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_B (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_D (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold104_X (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_SCD (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold129_X (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_SCE (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold158_X (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net581));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
