module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net608;
 wire net645;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net843;
 wire clknet_1_0__leaf_net843;
 wire clknet_1_1__leaf_net843;
 wire clknet_0_net916;
 wire clknet_1_0__leaf_net916;
 wire clknet_1_1__leaf_net916;
 wire clknet_0_net746;
 wire clknet_1_0__leaf_net746;
 wire clknet_1_1__leaf_net746;
 wire clknet_0_net747;
 wire clknet_1_0__leaf_net747;
 wire clknet_1_1__leaf_net747;
 wire clknet_0_net821;
 wire clknet_1_0__leaf_net821;
 wire clknet_1_1__leaf_net821;
 wire clknet_0_net542;
 wire clknet_1_0__leaf_net542;
 wire clknet_1_1__leaf_net542;
 wire clknet_0_net842;
 wire clknet_1_0__leaf_net842;
 wire clknet_1_1__leaf_net842;
 wire clknet_0_net841;
 wire clknet_1_0__leaf_net841;
 wire clknet_1_1__leaf_net841;
 wire clknet_0_net604;
 wire clknet_1_0__leaf_net604;
 wire clknet_1_1__leaf_net604;
 wire clknet_0_net742;
 wire clknet_1_0__leaf_net742;
 wire clknet_1_1__leaf_net742;
 wire clknet_0_net823;
 wire clknet_1_0__leaf_net823;
 wire clknet_1_1__leaf_net823;
 wire clknet_0_net822;
 wire clknet_1_0__leaf_net822;
 wire clknet_1_1__leaf_net822;
 wire clknet_0_net537;
 wire clknet_1_0__leaf_net537;
 wire clknet_1_1__leaf_net537;
 wire clknet_0_net805;
 wire clknet_1_0__leaf_net805;
 wire clknet_1_1__leaf_net805;
 wire clknet_0_net534;
 wire clknet_1_0__leaf_net534;
 wire clknet_1_1__leaf_net534;
 wire clknet_0_net485;
 wire clknet_1_0__leaf_net485;
 wire clknet_1_1__leaf_net485;
 wire clknet_0_net804;
 wire clknet_1_0__leaf_net804;
 wire clknet_1_1__leaf_net804;
 wire clknet_0_net618;
 wire clknet_1_0__leaf_net618;
 wire clknet_1_1__leaf_net618;
 wire clknet_0_net803;
 wire clknet_1_0__leaf_net803;
 wire clknet_1_1__leaf_net803;
 wire clknet_0_net498;
 wire clknet_1_0__leaf_net498;
 wire clknet_1_1__leaf_net498;
 wire clknet_0_net477;
 wire clknet_1_0__leaf_net477;
 wire clknet_1_1__leaf_net477;
 wire clknet_0_net581;
 wire clknet_1_0__leaf_net581;
 wire clknet_1_1__leaf_net581;
 wire clknet_0_net575;
 wire clknet_1_0__leaf_net575;
 wire clknet_1_1__leaf_net575;
 wire clknet_0_net568;
 wire clknet_1_0__leaf_net568;
 wire clknet_1_1__leaf_net568;
 wire clknet_0_net787;
 wire clknet_1_0__leaf_net787;
 wire clknet_1_1__leaf_net787;
 wire clknet_0_net380;
 wire clknet_1_0__leaf_net380;
 wire clknet_1_1__leaf_net380;
 wire clknet_0_net496;
 wire clknet_1_0__leaf_net496;
 wire clknet_1_1__leaf_net496;
 wire clknet_0_net479;
 wire clknet_1_0__leaf_net479;
 wire clknet_1_1__leaf_net479;
 wire clknet_0_net400;
 wire clknet_1_0__leaf_net400;
 wire clknet_1_1__leaf_net400;
 wire clknet_0_net507;
 wire clknet_1_0__leaf_net507;
 wire clknet_1_1__leaf_net507;
 wire clknet_0_net399;
 wire clknet_1_0__leaf_net399;
 wire clknet_1_1__leaf_net399;
 wire clknet_0_net372;
 wire clknet_1_0__leaf_net372;
 wire clknet_1_1__leaf_net372;
 wire clknet_0_net951;
 wire clknet_1_0__leaf_net951;
 wire clknet_1_1__leaf_net951;
 wire clknet_0_net361;
 wire clknet_1_0__leaf_net361;
 wire clknet_1_1__leaf_net361;
 wire clknet_0_net786;
 wire clknet_1_0__leaf_net786;
 wire clknet_1_1__leaf_net786;
 wire clknet_0_net569;
 wire clknet_1_0__leaf_net569;
 wire clknet_1_1__leaf_net569;
 wire clknet_0_net567;
 wire clknet_1_0__leaf_net567;
 wire clknet_1_1__leaf_net567;
 wire clknet_0_net768;
 wire clknet_1_0__leaf_net768;
 wire clknet_1_1__leaf_net768;
 wire clknet_0_net389;
 wire clknet_1_0__leaf_net389;
 wire clknet_1_1__leaf_net389;
 wire clknet_0_net269;
 wire clknet_1_0__leaf_net269;
 wire clknet_1_1__leaf_net269;
 wire clknet_0_net264;
 wire clknet_1_0__leaf_net264;
 wire clknet_1_1__leaf_net264;
 wire clknet_0_net254;
 wire clknet_1_0__leaf_net254;
 wire clknet_1_1__leaf_net254;
 wire clknet_0_net767;
 wire clknet_1_0__leaf_net767;
 wire clknet_1_1__leaf_net767;
 wire clknet_0_net396;
 wire clknet_1_0__leaf_net396;
 wire clknet_1_1__leaf_net396;
 wire clknet_0_net913;
 wire clknet_1_0__leaf_net913;
 wire clknet_1_1__leaf_net913;
 wire clknet_0_net378;
 wire clknet_1_0__leaf_net378;
 wire clknet_1_1__leaf_net378;
 wire clknet_0_net365;
 wire clknet_1_0__leaf_net365;
 wire clknet_1_1__leaf_net365;
 wire clknet_0_net275;
 wire clknet_1_0__leaf_net275;
 wire clknet_1_1__leaf_net275;
 wire clknet_0_net230;
 wire clknet_1_0__leaf_net230;
 wire clknet_1_1__leaf_net230;
 wire clknet_0_net706;
 wire clknet_1_0__leaf_net706;
 wire clknet_1_1__leaf_net706;
 wire clknet_0_net570;
 wire clknet_1_0__leaf_net570;
 wire clknet_1_1__leaf_net570;
 wire clknet_0_net392;
 wire clknet_1_0__leaf_net392;
 wire clknet_1_1__leaf_net392;
 wire clknet_0_net343;
 wire clknet_1_0__leaf_net343;
 wire clknet_1_1__leaf_net343;
 wire clknet_0_net366;
 wire clknet_1_0__leaf_net366;
 wire clknet_1_1__leaf_net366;
 wire clknet_0_net354;
 wire clknet_1_0__leaf_net354;
 wire clknet_1_1__leaf_net354;
 wire clknet_0_net349;
 wire clknet_1_0__leaf_net349;
 wire clknet_1_1__leaf_net349;
 wire clknet_0_net233;
 wire clknet_1_0__leaf_net233;
 wire clknet_1_1__leaf_net233;
 wire clknet_0_net232;
 wire clknet_1_0__leaf_net232;
 wire clknet_1_1__leaf_net232;
 wire clknet_0_net952;
 wire clknet_1_0__leaf_net952;
 wire clknet_1_1__leaf_net952;
 wire clknet_0_net280;
 wire clknet_1_0__leaf_net280;
 wire clknet_1_1__leaf_net280;
 wire clknet_0_net925;
 wire clknet_1_0__leaf_net925;
 wire clknet_1_1__leaf_net925;
 wire clknet_0_net953;
 wire clknet_1_0__leaf_net953;
 wire clknet_1_1__leaf_net953;
 wire clknet_0_net316;
 wire clknet_1_0__leaf_net316;
 wire clknet_1_1__leaf_net316;
 wire clknet_0_net948;
 wire clknet_1_0__leaf_net948;
 wire clknet_1_1__leaf_net948;
 wire clknet_0_net299;
 wire clknet_1_0__leaf_net299;
 wire clknet_1_1__leaf_net299;
 wire clknet_0_net308;
 wire clknet_1_0__leaf_net308;
 wire clknet_1_1__leaf_net308;
 wire clknet_0_net188;
 wire clknet_1_0__leaf_net188;
 wire clknet_1_1__leaf_net188;
 wire clknet_0_net189;
 wire clknet_1_0__leaf_net189;
 wire clknet_1_1__leaf_net189;
 wire clknet_0_net177;
 wire clknet_1_0__leaf_net177;
 wire clknet_1_1__leaf_net177;
 wire clknet_0_net178;
 wire clknet_1_0__leaf_net178;
 wire clknet_1_1__leaf_net178;
 wire clknet_0_net930;
 wire clknet_1_0__leaf_net930;
 wire clknet_1_1__leaf_net930;
 wire clknet_0_net182;
 wire clknet_1_0__leaf_net182;
 wire clknet_1_1__leaf_net182;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;

 sky130_fd_sc_hd__or4bb_1 c100 (.A(net26),
    .B(net34),
    .C_N(net29),
    .D_N(net6),
    .X(net38));
 sky130_fd_sc_hd__and3_4 c101 (.A(net30),
    .B(net27),
    .C(net1024),
    .X(net39));
 sky130_fd_sc_hd__or4bb_4 c102 (.A(net2),
    .B(net1032),
    .C_N(net1018),
    .D_N(net38),
    .X(net40));
 sky130_fd_sc_hd__a2111o_2 c103 (.A1(net35),
    .A2(net34),
    .B1(net38),
    .C1(net40),
    .D1(net27),
    .X(net41));
 sky130_fd_sc_hd__mux4_2 c104 (.A0(net39),
    .A1(net981),
    .A2(net34),
    .A3(net894),
    .S0(net37),
    .S1(net26),
    .X(net42));
 sky130_fd_sc_hd__mux4_2 c105 (.A0(net874),
    .A1(net41),
    .A2(net40),
    .A3(net13),
    .S0(net42),
    .S1(net36),
    .X(net939));
 sky130_fd_sc_hd__mux4_2 c106 (.A0(net37),
    .A1(net30),
    .A2(net40),
    .A3(net1029),
    .S0(net33),
    .S1(net41),
    .X(net43));
 sky130_fd_sc_hd__mux4_2 c107 (.A0(net29),
    .A1(net25),
    .A2(net39),
    .A3(net939),
    .S0(net36),
    .S1(net43),
    .X(net44));
 sky130_fd_sc_hd__mux4_2 c108 (.A0(net38),
    .A1(net887),
    .A2(net42),
    .A3(net44),
    .S0(net39),
    .S1(net31),
    .X(net45));
 sky130_fd_sc_hd__mux4_2 c109 (.A0(net45),
    .A1(net1085),
    .A2(net939),
    .A3(net27),
    .S0(net30),
    .S1(net44),
    .X(net46));
 sky130_fd_sc_hd__and3_1 c110 (.A(net30),
    .B(net1021),
    .C(net1028),
    .X(net47));
 sky130_fd_sc_hd__or4bb_1 c111 (.A(net15),
    .B(net47),
    .C_N(net882),
    .D_N(net25),
    .X(net48));
 sky130_fd_sc_hd__and3_1 c112 (.A(net882),
    .B(net1033),
    .C(net25),
    .X(net49));
 sky130_fd_sc_hd__and3_2 c113 (.A(net29),
    .B(net37),
    .C(net1032),
    .X(net50));
 sky130_fd_sc_hd__and3_1 c114 (.A(net35),
    .B(net48),
    .C(net1024),
    .X(net51));
 sky130_fd_sc_hd__and3_1 c115 (.A(net1040),
    .B(net49),
    .C(net1020),
    .X(net52));
 sky130_fd_sc_hd__a2111o_1 c116 (.A1(net51),
    .A2(net6),
    .B1(net32),
    .C1(net1021),
    .D1(net1024),
    .X(net53));
 sky130_fd_sc_hd__and3_1 c117 (.A(net52),
    .B(net15),
    .C(net50),
    .X(net54));
 sky130_fd_sc_hd__a2111o_4 c118 (.A1(net883),
    .A2(net10),
    .B1(net30),
    .C1(net1035),
    .D1(net36),
    .X(net55));
 sky130_fd_sc_hd__and3_1 c119 (.A(net49),
    .B(net1033),
    .C(net50),
    .X(net56));
 sky130_fd_sc_hd__and3_1 c120 (.A(net56),
    .B(net30),
    .C(net1130),
    .X(net57));
 sky130_fd_sc_hd__and3_2 c121 (.A(net1045),
    .B(net861),
    .C(net1026),
    .X(net943));
 sky130_fd_sc_hd__or4bb_1 c122 (.A(net865),
    .B(net41),
    .C_N(net883),
    .D_N(net57),
    .X(net58));
 sky130_fd_sc_hd__mux4_1 c123 (.A0(net47),
    .A1(net52),
    .A2(net939),
    .A3(net987),
    .S0(net56),
    .S1(net50),
    .X(net59));
 sky130_fd_sc_hd__a2111o_1 c124 (.A1(net59),
    .A2(net883),
    .B1(net51),
    .C1(net41),
    .D1(net1032),
    .X(net60));
 sky130_fd_sc_hd__a2111o_1 c125 (.A1(net41),
    .A2(net939),
    .B1(net59),
    .C1(net57),
    .D1(net1024),
    .X(net61));
 sky130_fd_sc_hd__and3_1 c126 (.A(net57),
    .B(net1033),
    .C(net1087),
    .X(net62));
 sky130_fd_sc_hd__a2111o_1 c127 (.A1(net60),
    .A2(net29),
    .B1(net58),
    .C1(net62),
    .D1(net54),
    .X(net63));
 sky130_fd_sc_hd__and3_4 c128 (.A(net54),
    .B(net55),
    .C(net943),
    .X(net64));
 sky130_fd_sc_hd__mux4_1 c129 (.A0(net62),
    .A1(net58),
    .A2(net1040),
    .A3(net50),
    .S0(net49),
    .S1(net943),
    .X(net65));
 sky130_fd_sc_hd__mux4_1 c130 (.A0(net63),
    .A1(net943),
    .A2(net64),
    .A3(net42),
    .S0(net1087),
    .S1(net65),
    .X(net66));
 sky130_fd_sc_hd__mux4_2 c131 (.A0(net65),
    .A1(net66),
    .A2(net64),
    .A3(net63),
    .S0(net1040),
    .S1(net60),
    .X(net67));
 sky130_fd_sc_hd__and3_1 c132 (.A(net1045),
    .B(net1046),
    .C(net1027),
    .X(net929));
 sky130_fd_sc_hd__and3_4 c133 (.A(net903),
    .B(net1041),
    .C(net1044),
    .X(net68));
 sky130_fd_sc_hd__and3_4 c134 (.A(net1040),
    .B(net1038),
    .C(net1027),
    .X(net69));
 sky130_fd_sc_hd__and2_4 c135 (.A(net904),
    .B(net1038),
    .X(net70));
 sky130_fd_sc_hd__and3_4 c136 (.A(net1013),
    .B(net1040),
    .C(net1023),
    .X(net71));
 sky130_fd_sc_hd__or4bb_1 c137 (.A(net1036),
    .B(net69),
    .C_N(net1046),
    .D_N(net1034),
    .X(net72));
 sky130_fd_sc_hd__and3_4 c138 (.A(net71),
    .B(net1027),
    .C(net1040),
    .X(net73));
 sky130_fd_sc_hd__and3_2 c139 (.A(net1013),
    .B(net858),
    .C(net1001),
    .X(net74));
 sky130_fd_sc_hd__or4bb_4 c140 (.A(net858),
    .B(net1038),
    .C_N(net1001),
    .D_N(net1013),
    .X(net75));
 sky130_fd_sc_hd__and3_4 c141 (.A(net73),
    .B(net1041),
    .C(net1002),
    .X(net76));
 sky130_fd_sc_hd__and3_4 c142 (.A(net997),
    .B(net1013),
    .C(net1043),
    .X(net77));
 sky130_fd_sc_hd__a2111o_1 c143 (.A1(net997),
    .A2(net1041),
    .B1(net1016),
    .C1(net1046),
    .D1(net1001),
    .X(net78));
 sky130_fd_sc_hd__and3_1 c144 (.A(net996),
    .B(net1046),
    .C(net997),
    .X(net910));
 sky130_fd_sc_hd__mux4_2 c145 (.A0(net71),
    .A1(net904),
    .A2(net992),
    .A3(net996),
    .S0(net1013),
    .S1(net1001),
    .X(net79));
 sky130_fd_sc_hd__and3_4 c146 (.A(net1106),
    .B(net1046),
    .C(net73),
    .X(net80));
 sky130_fd_sc_hd__mux4_2 c147 (.A0(net992),
    .A1(net75),
    .A2(net80),
    .A3(net73),
    .S0(net74),
    .S1(net1002),
    .X(net81));
 sky130_fd_sc_hd__or4bb_4 c148 (.A(net997),
    .B(net990),
    .C_N(net1034),
    .D_N(net1001),
    .X(net82));
 sky130_fd_sc_hd__and3_2 c149 (.A(net74),
    .B(net68),
    .C(net1106),
    .X(net83));
 sky130_fd_sc_hd__or4bb_4 c150 (.A(net1106),
    .B(net71),
    .C_N(net1018),
    .D_N(net990),
    .X(net84));
 sky130_fd_sc_hd__a2111o_4 c151 (.A1(net1001),
    .A2(net74),
    .B1(net83),
    .C1(net1046),
    .D1(net1106),
    .X(net85));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net989),
    .A1(net83),
    .A2(net85),
    .A3(net1001),
    .S0(net69),
    .S1(net1013),
    .X(net86));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net86),
    .A1(net990),
    .A2(net75),
    .A3(net80),
    .S0(net79),
    .S1(net1013),
    .X(net87));
 sky130_fd_sc_hd__or4bb_1 c154 (.A(net1037),
    .B(net864),
    .C_N(net872),
    .D_N(net869),
    .X(net932));
 sky130_fd_sc_hd__a2111o_1 c155 (.A1(net876),
    .A2(net1034),
    .B1(net882),
    .C1(net1002),
    .D1(net1038),
    .X(net88));
 sky130_fd_sc_hd__and3_1 c156 (.A(net871),
    .B(net83),
    .C(net877),
    .X(net89));
 sky130_fd_sc_hd__mux4_2 c157 (.A0(net880),
    .A1(net1027),
    .A2(net1013),
    .A3(net71),
    .S0(net870),
    .S1(net1011),
    .X(net90));
 sky130_fd_sc_hd__and3_1 c158 (.A(net90),
    .B(net872),
    .C(net86),
    .X(net91));
 sky130_fd_sc_hd__and3_1 c159 (.A(net1041),
    .B(net90),
    .C(net873),
    .X(net92));
 sky130_fd_sc_hd__and3_2 c160 (.A(net89),
    .B(net92),
    .C(net870),
    .X(net93));
 sky130_fd_sc_hd__mux4_2 c161 (.A0(net92),
    .A1(net86),
    .A2(net69),
    .A3(net990),
    .S0(net1011),
    .S1(net1045),
    .X(net94));
 sky130_fd_sc_hd__mux4_2 c162 (.A0(net872),
    .A1(net94),
    .A2(net879),
    .A3(net1037),
    .S0(net881),
    .S1(net1011),
    .X(net95));
 sky130_fd_sc_hd__or4bb_4 c163 (.A(net1105),
    .B(net85),
    .C_N(net1106),
    .D_N(net1104),
    .X(net96));
 sky130_fd_sc_hd__or4bb_2 c164 (.A(net94),
    .B(net996),
    .C_N(net998),
    .D_N(net1002),
    .X(net97));
 sky130_fd_sc_hd__mux4_2 c165 (.A0(net853),
    .A1(net876),
    .A2(net96),
    .A3(net1011),
    .S0(net859),
    .S1(net94),
    .X(net98));
 sky130_fd_sc_hd__a2111o_1 c166 (.A1(net93),
    .A2(net862),
    .B1(net92),
    .C1(net1103),
    .D1(net1001),
    .X(net99));
 sky130_fd_sc_hd__a2111o_1 c167 (.A1(net1022),
    .A2(net866),
    .B1(net989),
    .C1(net1103),
    .D1(net94),
    .X(net100));
 sky130_fd_sc_hd__mux4_2 c168 (.A0(net998),
    .A1(net1042),
    .A2(net97),
    .A3(net69),
    .S0(net979),
    .S1(net984),
    .X(net101));
 sky130_fd_sc_hd__and3_1 c169 (.A(net1103),
    .B(net96),
    .C(net99),
    .X(net102));
 sky130_fd_sc_hd__mux4_2 c170 (.A0(net101),
    .A1(net85),
    .A2(net877),
    .A3(net865),
    .S0(net1103),
    .S1(net80),
    .X(net103));
 sky130_fd_sc_hd__a2111o_4 c171 (.A1(net103),
    .A2(net862),
    .B1(net871),
    .C1(net1103),
    .D1(net101),
    .X(net104));
 sky130_fd_sc_hd__mux4_2 c172 (.A0(net99),
    .A1(net104),
    .A2(net89),
    .A3(net102),
    .S0(net101),
    .S1(net103),
    .X(net105));
 sky130_fd_sc_hd__or4bb_4 c173 (.A(net104),
    .B(net99),
    .C_N(net100),
    .D_N(net1103),
    .X(net106));
 sky130_fd_sc_hd__and3_4 c174 (.A(net974),
    .B(net100),
    .C(net1103),
    .X(net107));
 sky130_fd_sc_hd__mux4_2 c175 (.A0(net107),
    .A1(net1065),
    .A2(net974),
    .A3(net872),
    .S0(net873),
    .S1(net979),
    .X(net108));
 sky130_fd_sc_hd__or4bb_2 c176 (.A(net100),
    .B(net881),
    .C_N(net902),
    .D_N(net1025),
    .X(net109));
 sky130_fd_sc_hd__or4bb_4 c177 (.A(net0),
    .B(net896),
    .C_N(net101),
    .D_N(net974),
    .X(net110));
 sky130_fd_sc_hd__a2111o_4 c178 (.A1(net881),
    .A2(net1029),
    .B1(net888),
    .C1(net1106),
    .D1(net901),
    .X(net111));
 sky130_fd_sc_hd__and3_1 c179 (.A(net89),
    .B(net1124),
    .C(net899),
    .X(net112));
 sky130_fd_sc_hd__and3_1 c180 (.A(net99),
    .B(net111),
    .C(net105),
    .X(net113));
 sky130_fd_sc_hd__and3_4 c181 (.A(net90),
    .B(net989),
    .C(net111),
    .X(net114));
 sky130_fd_sc_hd__a2111o_4 c182 (.A1(net872),
    .A2(net114),
    .B1(net110),
    .C1(net1061),
    .D1(net1090),
    .X(net115));
 sky130_fd_sc_hd__or4bb_4 c183 (.A(net113),
    .B(net1124),
    .C_N(net111),
    .D_N(net871),
    .X(net116));
 sky130_fd_sc_hd__or4bb_4 c184 (.A(net872),
    .B(net112),
    .C_N(net968),
    .D_N(net1065),
    .X(net117));
 sky130_fd_sc_hd__and3_2 c185 (.A(net1036),
    .B(net1026),
    .C(net104),
    .X(net118));
 sky130_fd_sc_hd__or4bb_4 c186 (.A(net93),
    .B(net995),
    .C_N(net110),
    .D_N(net997),
    .X(net931));
 sky130_fd_sc_hd__or4bb_4 c187 (.A(net877),
    .B(net902),
    .C_N(net1011),
    .D_N(net118),
    .X(net119));
 sky130_fd_sc_hd__or4bb_2 c188 (.A(net119),
    .B(net116),
    .C_N(net94),
    .D_N(net113),
    .X(net120));
 sky130_fd_sc_hd__mux4_2 c189 (.A0(net83),
    .A1(net80),
    .A2(net896),
    .A3(net112),
    .S0(net967),
    .S1(net1025),
    .X(net121));
 sky130_fd_sc_hd__or4bb_2 c190 (.A(net101),
    .B(net120),
    .C_N(net904),
    .D_N(net118),
    .X(net122));
 sky130_fd_sc_hd__mux4_1 c191 (.A0(net117),
    .A1(net974),
    .A2(net122),
    .A3(net109),
    .S0(net1011),
    .S1(net115),
    .X(net123));
 sky130_fd_sc_hd__mux4_1 c192 (.A0(net118),
    .A1(net109),
    .A2(net120),
    .A3(net1017),
    .S0(net989),
    .S1(net122),
    .X(net124));
 sky130_fd_sc_hd__a2111o_2 c193 (.A1(net880),
    .A2(net102),
    .B1(net121),
    .C1(net99),
    .D1(net898),
    .X(net125));
 sky130_fd_sc_hd__a2111o_1 c194 (.A1(net122),
    .A2(net110),
    .B1(net120),
    .C1(net125),
    .D1(net116),
    .X(net126));
 sky130_fd_sc_hd__mux4_1 c195 (.A0(net898),
    .A1(net125),
    .A2(net112),
    .A3(net1038),
    .S0(net118),
    .S1(net685),
    .X(net127));
 sky130_fd_sc_hd__a2111o_1 c196 (.A1(net121),
    .A2(net979),
    .B1(net125),
    .C1(net686),
    .D1(net763),
    .X(net128));
 sky130_fd_sc_hd__mux4_2 c197 (.A0(net1057),
    .A1(net115),
    .A2(net114),
    .A3(net82),
    .S0(net686),
    .S1(net762),
    .X(net129));
 sky130_fd_sc_hd__or4bb_2 c198 (.A(net1124),
    .B(net112),
    .C_N(net998),
    .D_N(net866),
    .X(net130));
 sky130_fd_sc_hd__mux4_2 c199 (.A0(net22),
    .A1(net83),
    .A2(net989),
    .A3(net1076),
    .S0(net71),
    .S1(net1103),
    .X(net131));
 sky130_fd_sc_hd__a2111o_1 c200 (.A1(net80),
    .A2(net870),
    .B1(net120),
    .C1(net876),
    .D1(net974),
    .X(net132));
 sky130_fd_sc_hd__a2111o_1 c201 (.A1(net1086),
    .A2(net1033),
    .B1(net993),
    .C1(net1089),
    .D1(net682),
    .X(net133));
 sky130_fd_sc_hd__mux4_2 c202 (.A0(net11),
    .A1(net1034),
    .A2(net1035),
    .A3(net19),
    .S0(net997),
    .S1(net1014),
    .X(net134));
 sky130_fd_sc_hd__a2111o_1 c203 (.A1(net1016),
    .A2(net18),
    .B1(net1028),
    .C1(net20),
    .D1(net685),
    .X(net135));
 sky130_fd_sc_hd__a2111o_2 c204 (.A1(net9),
    .A2(net112),
    .B1(net16),
    .C1(net130),
    .D1(net993),
    .X(net136));
 sky130_fd_sc_hd__a2111o_2 c205 (.A1(net120),
    .A2(net133),
    .B1(net1104),
    .C1(net68),
    .D1(net1089),
    .X(net137));
 sky130_fd_sc_hd__mux4_1 c206 (.A0(net102),
    .A1(net134),
    .A2(net136),
    .A3(net901),
    .S0(net1106),
    .S1(net681),
    .X(net138));
 sky130_fd_sc_hd__sdfbbn_2 c207 (.CLK_N(clknet_4_2_0_clk),
    .D(net112),
    .RESET_B(net137),
    .SCD(net104),
    .SCE(net129),
    .SET_B(net14),
    .Q(net140),
    .Q_N(net139));
 sky130_fd_sc_hd__mux4_2 c208 (.A0(net135),
    .A1(net138),
    .A2(net6),
    .A3(net139),
    .S0(net70),
    .S1(net681),
    .X(net946));
 sky130_fd_sc_hd__a2111o_1 c209 (.A1(net997),
    .A2(net998),
    .B1(net138),
    .C1(net139),
    .D1(net82),
    .X(net141));
 sky130_fd_sc_hd__a2111o_1 c210 (.A1(net1010),
    .A2(net129),
    .B1(net137),
    .C1(net133),
    .D1(net1026),
    .X(net142));
 sky130_fd_sc_hd__a2111o_1 c211 (.A1(net83),
    .A2(net132),
    .B1(net1010),
    .C1(net1103),
    .D1(net1009),
    .X(net143));
 sky130_fd_sc_hd__a2111o_1 c212 (.A1(net869),
    .A2(net135),
    .B1(net107),
    .C1(net139),
    .D1(net664),
    .X(net144));
 sky130_fd_sc_hd__mux4_1 c213 (.A0(net141),
    .A1(net1121),
    .A2(net137),
    .A3(net1010),
    .S0(net16),
    .S1(net144),
    .X(net145));
 sky130_fd_sc_hd__mux4_2 c214 (.A0(net144),
    .A1(net136),
    .A2(net117),
    .A3(net102),
    .S0(net139),
    .S1(net763),
    .X(net146));
 sky130_fd_sc_hd__mux4_2 c215 (.A0(net138),
    .A1(net135),
    .A2(net131),
    .A3(net115),
    .S0(net664),
    .S1(net681),
    .X(net147));
 sky130_fd_sc_hd__mux4_1 c216 (.A0(net121),
    .A1(net133),
    .A2(net130),
    .A3(net147),
    .S0(net664),
    .S1(net1009),
    .X(net148));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(net148),
    .A1(net1010),
    .A2(net147),
    .A3(net146),
    .S0(net1104),
    .S1(net979),
    .X(net149));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(net136),
    .A1(net138),
    .A2(net6),
    .A3(net148),
    .S0(net681),
    .S1(net1009),
    .X(net150));
 sky130_fd_sc_hd__a2111o_1 c219 (.A1(net144),
    .A2(net131),
    .B1(net115),
    .C1(net664),
    .D1(net1009),
    .X(net151));
 sky130_fd_sc_hd__a2111o_4 c220 (.A1(net901),
    .A2(net1073),
    .B1(net1029),
    .C1(net1023),
    .D1(net1016),
    .X(net908));
 sky130_fd_sc_hd__a2111o_4 c221 (.A1(net151),
    .A2(net111),
    .B1(net1128),
    .C1(net887),
    .D1(net901),
    .X(net927));
 sky130_fd_sc_hd__a2111o_1 c222 (.A1(net129),
    .A2(net1104),
    .B1(net40),
    .C1(net1025),
    .D1(net1103),
    .X(net152));
 sky130_fd_sc_hd__a2111o_1 c223 (.A1(net40),
    .A2(net80),
    .B1(net1010),
    .C1(net1077),
    .D1(net1014),
    .X(net153));
 sky130_fd_sc_hd__mux4_1 c224 (.A0(net903),
    .A1(net1079),
    .A2(net991),
    .A3(net893),
    .S0(net1001),
    .S1(net139),
    .X(net154));
 sky130_fd_sc_hd__mux4_2 c225 (.A0(net154),
    .A1(net967),
    .A2(net1010),
    .A3(net4),
    .S0(net1032),
    .S1(net1043),
    .X(net155));
 sky130_fd_sc_hd__a2111o_1 c226 (.A1(net155),
    .A2(net33),
    .B1(net968),
    .C1(net927),
    .D1(net908),
    .X(net156));
 sky130_fd_sc_hd__mux4_1 c227 (.A0(net111),
    .A1(net155),
    .A2(net151),
    .A3(net989),
    .S0(net927),
    .S1(net664),
    .X(net157));
 sky130_fd_sc_hd__a2111o_1 c228 (.A1(net152),
    .A2(net151),
    .B1(net927),
    .C1(net1042),
    .D1(net1033),
    .X(net158));
 sky130_fd_sc_hd__a2111o_1 c229 (.A1(net16),
    .A2(net1084),
    .B1(net1),
    .C1(net1076),
    .D1(net927),
    .X(net159));
 sky130_fd_sc_hd__mux4_1 c230 (.A0(net155),
    .A1(net1023),
    .A2(net1042),
    .A3(net43),
    .S0(net152),
    .S1(net663),
    .X(net160));
 sky130_fd_sc_hd__a2111o_1 c231 (.A1(net146),
    .A2(net1084),
    .B1(net1107),
    .C1(net663),
    .D1(net761),
    .X(net161));
 sky130_fd_sc_hd__mux4_1 c232 (.A0(net7),
    .A1(net155),
    .A2(net1085),
    .A3(net1080),
    .S0(net154),
    .S1(net692),
    .X(net162));
 sky130_fd_sc_hd__sdfbbn_2 c233 (.CLK_N(clknet_4_0_0_clk),
    .D(net1130),
    .RESET_B(net46),
    .SCD(net152),
    .SCE(net663),
    .SET_B(net664),
    .Q(net933),
    .Q_N(net163));
 sky130_fd_sc_hd__mux4_1 c234 (.A0(net1080),
    .A1(net1059),
    .A2(net1010),
    .A3(net1032),
    .S0(net692),
    .S1(net761),
    .X(net164));
 sky130_fd_sc_hd__mux4_1 c235 (.A0(net164),
    .A1(net0),
    .A2(net162),
    .A3(net908),
    .S0(net111),
    .S1(net718),
    .X(net165));
 sky130_fd_sc_hd__a2111o_1 c236 (.A1(net115),
    .A2(net163),
    .B1(net974),
    .C1(net718),
    .D1(net752),
    .X(net166));
 sky130_fd_sc_hd__mux4_1 c237 (.A0(net1060),
    .A1(net146),
    .A2(net166),
    .A3(net162),
    .S0(net718),
    .S1(net761),
    .X(net167));
 sky130_fd_sc_hd__mux4_1 c238 (.A0(net80),
    .A1(net10),
    .A2(net129),
    .A3(net927),
    .S0(net139),
    .S1(net765),
    .X(net168));
 sky130_fd_sc_hd__mux4_2 c239 (.A0(net43),
    .A1(net153),
    .A2(net114),
    .A3(net33),
    .S0(net765),
    .S1(net766),
    .X(net169));
 sky130_fd_sc_hd__mux4_2 c240 (.A0(net129),
    .A1(net131),
    .A2(net1070),
    .A3(net968),
    .S0(net663),
    .S1(net762),
    .X(net170));
 sky130_fd_sc_hd__sdfbbp_1 c241 (.CLK(clknet_4_1_0_clk),
    .D(net166),
    .RESET_B(net170),
    .SCD(net164),
    .SCE(net1033),
    .SET_B(net1093),
    .Q(net172),
    .Q_N(net171));
 sky130_fd_sc_hd__mux4_1 c242 (.A0(clknet_1_0__leaf_net188),
    .A1(net48),
    .A2(net943),
    .A3(clknet_1_0__leaf_net189),
    .S0(net1024),
    .S1(net766),
    .X(net173));
 sky130_fd_sc_hd__mux4_2 c243 (.A0(net25),
    .A1(net36),
    .A2(net939),
    .A3(net1012),
    .S0(net1021),
    .S1(net1009),
    .X(net914));
 sky130_fd_sc_hd__mux4_1 c244 (.A0(net162),
    .A1(clknet_1_1__leaf_net188),
    .A2(net36),
    .A3(net1045),
    .S0(net1085),
    .S1(net190),
    .X(net174));
 sky130_fd_sc_hd__mux4_1 c245 (.A0(clknet_1_1__leaf_net189),
    .A1(net1024),
    .A2(net927),
    .A3(net914),
    .S0(net1051),
    .S1(net1014),
    .X(net175));
 sky130_fd_sc_hd__mux4_2 c246 (.A0(net1051),
    .A1(net0),
    .A2(net1014),
    .A3(net942),
    .S0(net674),
    .S1(net692),
    .X(net176));
 sky130_fd_sc_hd__mux4_1 c247 (.A0(net48),
    .A1(net1018),
    .A2(net674),
    .A3(net1009),
    .S0(net692),
    .S1(clknet_1_0__leaf_net925),
    .X(net177));
 sky130_fd_sc_hd__mux4_2 c248 (.A0(net176),
    .A1(clknet_1_1__leaf_net177),
    .A2(net55),
    .A3(net981),
    .S0(net673),
    .S1(net766),
    .X(net178));
 sky130_fd_sc_hd__mux4_1 c249 (.A0(net191),
    .A1(net860),
    .A2(net1087),
    .A3(net943),
    .S0(net1035),
    .S1(net765),
    .X(net179));
 sky130_fd_sc_hd__mux4_1 c250 (.A0(net131),
    .A1(net179),
    .A2(net967),
    .A3(net53),
    .S0(net1018),
    .S1(net1040),
    .X(net180));
 sky130_fd_sc_hd__mux4_2 c251 (.A0(net1035),
    .A1(net55),
    .A2(net1085),
    .A3(net53),
    .S0(net699),
    .S1(net765),
    .X(net181));
 sky130_fd_sc_hd__mux4_1 c252 (.A0(net1087),
    .A1(net914),
    .A2(net176),
    .A3(clknet_1_0__leaf_net178),
    .S0(net55),
    .S1(net987),
    .X(net930));
 sky130_fd_sc_hd__mux4_1 c253 (.A0(net191),
    .A1(net36),
    .A2(clknet_1_0__leaf_net930),
    .A3(net163),
    .S0(net1088),
    .S1(net673),
    .X(net182));
 sky130_fd_sc_hd__mux4_1 c254 (.A0(clknet_1_1__leaf_net178),
    .A1(clknet_1_0__leaf_net182),
    .A2(clknet_1_1__leaf_net930),
    .A3(net1026),
    .S1(clknet_1_1__leaf_net925),
    .X(net183));
 sky130_fd_sc_hd__mux4_1 c255 (.A0(net10),
    .A1(clknet_1_0__leaf_net177),
    .A2(net186),
    .A3(net53),
    .S0(net170),
    .S1(net914),
    .X(net184));
 sky130_fd_sc_hd__mux4_1 c256 (.A0(net48),
    .A1(clknet_1_1__leaf_net188),
    .A2(net176),
    .A3(net1077),
    .S0(clknet_1_0__leaf_net182),
    .S1(net940),
    .X(net185));
 sky130_fd_sc_hd__mux4_1 c257 (.A0(net36),
    .A1(net1024),
    .A2(net1087),
    .A3(net865),
    .S0(net1077),
    .S1(net1021),
    .X(net186));
 sky130_fd_sc_hd__mux4_2 c258 (.A0(net53),
    .A1(net882),
    .A2(net64),
    .A3(net1024),
    .S0(net987),
    .S1(net1018),
    .X(net942));
 sky130_fd_sc_hd__mux4_1 c259 (.A0(net115),
    .A1(net861),
    .A2(net1032),
    .A3(net170),
    .S0(net1045),
    .S1(net1014),
    .X(net187));
 sky130_fd_sc_hd__mux4_1 c260 (.A0(net64),
    .A1(net67),
    .A2(net1014),
    .A3(net1077),
    .S0(net1035),
    .S1(clknet_1_0__leaf_net925),
    .X(net188));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(clknet_1_0__leaf_net188),
    .A1(net865),
    .A2(net993),
    .A3(net64),
    .S0(net115),
    .S1(net1009),
    .X(net189));
 sky130_fd_sc_hd__mux4_1 c262 (.A0(net186),
    .A1(net865),
    .A2(net1033),
    .A3(net64),
    .S0(net1077),
    .S1(net765),
    .X(net190));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net190),
    .A1(net1014),
    .A2(net1130),
    .A3(net1032),
    .S0(net1020),
    .S1(net967),
    .X(net191));
 sky130_fd_sc_hd__and3_1 c264 (.A(net903),
    .B(net1001),
    .C(net82),
    .X(net192));
 sky130_fd_sc_hd__and3_2 c265 (.A(net1043),
    .B(net74),
    .C(net192),
    .X(net193));
 sky130_fd_sc_hd__and3_4 c266 (.A(net1040),
    .B(net1018),
    .C(net1022),
    .X(net194));
 sky130_fd_sc_hd__and2_1 c267 (.A(net1039),
    .B(net1046),
    .X(net195));
 sky130_fd_sc_hd__mux4_2 c268 (.A0(net193),
    .A1(net1038),
    .A2(net990),
    .A3(net1043),
    .S0(net903),
    .S1(net1106),
    .X(net196));
 sky130_fd_sc_hd__and3_4 c269 (.A(net1034),
    .B(net192),
    .C(net77),
    .X(net197));
 sky130_fd_sc_hd__and3_2 c270 (.A(net193),
    .B(net195),
    .C(net996),
    .X(net198));
 sky130_fd_sc_hd__and2_2 c271 (.A(net193),
    .B(net75),
    .X(net199));
 sky130_fd_sc_hd__and3_1 c272 (.A(net199),
    .B(net196),
    .C(net1090),
    .X(net200));
 sky130_fd_sc_hd__and3_2 c273 (.A(net847),
    .B(net1039),
    .C(net199),
    .X(net201));
 sky130_fd_sc_hd__or4bb_4 c274 (.A(net192),
    .B(net1015),
    .C_N(net1016),
    .D_N(net1003),
    .X(net202));
 sky130_fd_sc_hd__and3_2 c275 (.A(net1046),
    .B(net79),
    .C(net193),
    .X(net203));
 sky130_fd_sc_hd__and3_4 c276 (.A(net201),
    .B(net202),
    .C(net200),
    .X(net204));
 sky130_fd_sc_hd__and3_2 c277 (.A(net197),
    .B(net201),
    .C(net193),
    .X(net205));
 sky130_fd_sc_hd__and3_2 c278 (.A(net205),
    .B(net199),
    .C(net203),
    .X(net206));
 sky130_fd_sc_hd__and3_1 c279 (.A(net858),
    .B(net205),
    .C(net202),
    .X(net207));
 sky130_fd_sc_hd__and3_1 c280 (.A(net206),
    .B(net207),
    .C(net1043),
    .X(net208));
 sky130_fd_sc_hd__and3_2 c281 (.A(net200),
    .B(net1106),
    .C(net975),
    .X(net209));
 sky130_fd_sc_hd__and3_1 c282 (.A(net209),
    .B(net206),
    .C(net975),
    .X(net210));
 sky130_fd_sc_hd__mux4_2 c283 (.A0(net1031),
    .A1(net207),
    .A2(net209),
    .A3(net975),
    .S0(net206),
    .S1(net194),
    .X(net211));
 sky130_fd_sc_hd__and3_2 c284 (.A(net198),
    .B(net211),
    .C(net972),
    .X(net212));
 sky130_fd_sc_hd__and3_4 c285 (.A(net212),
    .B(net203),
    .C(net211),
    .X(net213));
 sky130_fd_sc_hd__a2111o_1 c286 (.A1(net206),
    .A2(net103),
    .B1(net972),
    .C1(net1037),
    .D1(net1038),
    .X(net936));
 sky130_fd_sc_hd__and3_2 c287 (.A(net92),
    .B(net873),
    .C(net199),
    .X(net214));
 sky130_fd_sc_hd__or4bb_2 c288 (.A(net1015),
    .B(net992),
    .C_N(net980),
    .D_N(net969),
    .X(net215));
 sky130_fd_sc_hd__or4bb_4 c289 (.A(net989),
    .B(net92),
    .C_N(net969),
    .D_N(net200),
    .X(net216));
 sky130_fd_sc_hd__mux4_1 c290 (.A0(net1017),
    .A1(net201),
    .A2(net216),
    .A3(net108),
    .S0(net203),
    .S1(net969),
    .X(net217));
 sky130_fd_sc_hd__a2111o_2 c291 (.A1(net864),
    .A2(net1017),
    .B1(net1104),
    .C1(net107),
    .D1(net969),
    .X(net218));
 sky130_fd_sc_hd__and3_2 c292 (.A(net861),
    .B(net87),
    .C(net1002),
    .X(net219));
 sky130_fd_sc_hd__or4bb_2 c293 (.A(net214),
    .B(net873),
    .C_N(net992),
    .D_N(net969),
    .X(net220));
 sky130_fd_sc_hd__a2111o_4 c294 (.A1(net201),
    .A2(net998),
    .B1(net215),
    .C1(net992),
    .D1(net69),
    .X(net221));
 sky130_fd_sc_hd__mux4_2 c295 (.A0(net79),
    .A1(net93),
    .A2(net1046),
    .A3(net214),
    .S0(net216),
    .S1(net1037),
    .X(net222));
 sky130_fd_sc_hd__a2111o_1 c296 (.A1(net221),
    .A2(net217),
    .B1(net203),
    .C1(net103),
    .D1(net214),
    .X(net223));
 sky130_fd_sc_hd__and3_1 c297 (.A(net222),
    .B(net107),
    .C(net108),
    .X(net224));
 sky130_fd_sc_hd__a2111o_2 c298 (.A1(net217),
    .A2(net214),
    .B1(net88),
    .C1(net969),
    .D1(net979),
    .X(net957));
 sky130_fd_sc_hd__mux4_1 c299 (.A0(net85),
    .A1(net969),
    .A2(net972),
    .A3(net201),
    .S0(net220),
    .S1(net965),
    .X(net225));
 sky130_fd_sc_hd__a2111o_1 c300 (.A1(net870),
    .A2(net965),
    .B1(net863),
    .C1(net223),
    .D1(net214),
    .X(net226));
 sky130_fd_sc_hd__sdfrbp_2 c301 (.CLK(clknet_4_8_0_clk),
    .D(net1112),
    .RESET_B(net219),
    .SCD(net965),
    .SCE(clknet_1_1__leaf_net767),
    .Q(net918),
    .Q_N(net227));
 sky130_fd_sc_hd__or4bb_1 c302 (.A(net873),
    .B(net222),
    .C_N(net223),
    .D_N(net969),
    .X(net228));
 sky130_fd_sc_hd__mux4_1 c303 (.A0(net220),
    .A1(net196),
    .A2(net219),
    .A3(net200),
    .S0(net1062),
    .S1(net965),
    .X(net229));
 sky130_fd_sc_hd__a2111o_1 c304 (.A1(net918),
    .A2(net1046),
    .B1(net1091),
    .C1(net1006),
    .D1(clknet_1_1__leaf_net767),
    .X(net230));
 sky130_fd_sc_hd__mux4_1 c305 (.A0(net223),
    .A1(net196),
    .A2(clknet_1_0__leaf_net230),
    .A3(net193),
    .S0(net990),
    .S1(net1006),
    .X(net231));
 sky130_fd_sc_hd__mux4_1 c306 (.A0(net102),
    .A1(clknet_1_0__leaf_net230),
    .A2(net206),
    .A3(net218),
    .S0(net1040),
    .S1(net1008),
    .X(net232));
 sky130_fd_sc_hd__mux4_1 c307 (.A0(net216),
    .A1(clknet_1_1__leaf_net232),
    .A2(net1047),
    .A3(net1035),
    .S0(clknet_1_0__leaf_net230),
    .S1(net1006),
    .X(net233));
 sky130_fd_sc_hd__a2111o_2 c308 (.A1(net204),
    .A2(net860),
    .B1(net97),
    .C1(net984),
    .D1(net1029),
    .X(net234));
 sky130_fd_sc_hd__sdfbbn_2 c309 (.CLK_N(clknet_4_9_0_clk),
    .D(net223),
    .RESET_B(net125),
    .SCD(net113),
    .SCE(net209),
    .SET_B(net1002),
    .Q(net921),
    .Q_N(net235));
 sky130_fd_sc_hd__sdfbbn_2 c310 (.CLK_N(clknet_4_3_0_clk),
    .D(net879),
    .RESET_B(net897),
    .SCD(net216),
    .SCE(net1091),
    .SET_B(clknet_1_0__leaf_net233),
    .Q(net237),
    .Q_N(net236));
 sky130_fd_sc_hd__a2111o_2 c311 (.A1(net217),
    .A2(net218),
    .B1(net1011),
    .C1(net117),
    .D1(net116),
    .X(net238));
 sky130_fd_sc_hd__sdfbbp_1 c312 (.CLK(clknet_4_9_0_clk),
    .D(net113),
    .RESET_B(net204),
    .SCD(net125),
    .SCE(net980),
    .SET_B(net970),
    .Q(net240),
    .Q_N(net239));
 sky130_fd_sc_hd__a2111o_4 c313 (.A1(net240),
    .A2(net85),
    .B1(net107),
    .C1(net972),
    .D1(net995),
    .X(net241));
 sky130_fd_sc_hd__a2111o_2 c314 (.A1(net97),
    .A2(net1032),
    .B1(net236),
    .C1(net96),
    .D1(net686),
    .X(net937));
 sky130_fd_sc_hd__a2111o_1 c315 (.A1(net122),
    .A2(net891),
    .B1(net1026),
    .C1(net998),
    .D1(net218),
    .X(net242));
 sky130_fd_sc_hd__a2111o_1 c316 (.A1(net109),
    .A2(net237),
    .B1(net88),
    .C1(net975),
    .D1(net235),
    .X(net243));
 sky130_fd_sc_hd__a2111o_4 c317 (.A1(net896),
    .A2(net241),
    .B1(net243),
    .C1(net70),
    .D1(net859),
    .X(net244));
 sky130_fd_sc_hd__a2111o_2 c318 (.A1(net118),
    .A2(net110),
    .B1(net239),
    .C1(net234),
    .D1(net241),
    .X(net245));
 sky130_fd_sc_hd__a2111o_4 c319 (.A1(net1038),
    .A2(net118),
    .B1(net977),
    .C1(net921),
    .D1(net114),
    .X(net246));
 sky130_fd_sc_hd__a2111o_1 c320 (.A1(net1026),
    .A2(net121),
    .B1(net216),
    .C1(net109),
    .D1(net884),
    .X(net247));
 sky130_fd_sc_hd__mux4_2 c321 (.A0(net237),
    .A1(net96),
    .A2(net1017),
    .A3(net244),
    .S0(net235),
    .S1(net1026),
    .X(net248));
 sky130_fd_sc_hd__mux4_1 c322 (.A0(net238),
    .A1(net247),
    .A2(net975),
    .A3(net110),
    .S0(net246),
    .S1(net1038),
    .X(net249));
 sky130_fd_sc_hd__a2111o_1 c323 (.A1(net1),
    .A2(net248),
    .B1(net119),
    .C1(net245),
    .D1(net866),
    .X(net250));
 sky130_fd_sc_hd__mux4_1 c324 (.A0(net125),
    .A1(net238),
    .A2(net1002),
    .A3(net886),
    .S0(net995),
    .S1(net1006),
    .X(net251));
 sky130_fd_sc_hd__mux4_1 c325 (.A0(net1013),
    .A1(net194),
    .A2(net921),
    .A3(net977),
    .S0(net246),
    .S1(net239),
    .X(net252));
 sky130_fd_sc_hd__a2111o_1 c326 (.A1(net252),
    .A2(net121),
    .B1(net236),
    .C1(net887),
    .D1(net997),
    .X(net253));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(net977),
    .A1(net252),
    .A2(net216),
    .A3(net245),
    .S0(net1006),
    .S1(clknet_1_0__leaf_net768),
    .X(net254));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(net884),
    .A1(net246),
    .A2(net252),
    .A3(net1038),
    .S0(net235),
    .S1(net712),
    .X(net255));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net255),
    .A1(net247),
    .A2(net253),
    .A3(clknet_1_1__leaf_net254),
    .S0(net224),
    .S1(clknet_1_0__leaf_net767),
    .X(net256));
 sky130_fd_sc_hd__mux4_1 c330 (.A0(net133),
    .A1(net141),
    .A2(net93),
    .A3(net68),
    .S0(clknet_1_0__leaf_net254),
    .S1(net1004),
    .X(net257));
 sky130_fd_sc_hd__mux4_2 c331 (.A0(net998),
    .A1(net968),
    .A2(net921),
    .A3(net997),
    .S0(net8),
    .S1(net139),
    .X(net258));
 sky130_fd_sc_hd__mux4_1 c332 (.A0(net4),
    .A1(clknet_1_0__leaf_net232),
    .A2(net998),
    .A3(net227),
    .S0(net132),
    .S1(net949),
    .X(net259));
 sky130_fd_sc_hd__mux4_1 c333 (.A0(net245),
    .A1(clknet_1_0__leaf_net254),
    .A2(net235),
    .A3(net903),
    .S0(net234),
    .S1(clknet_1_0__leaf_net767),
    .X(net260));
 sky130_fd_sc_hd__mux4_1 c334 (.A0(net199),
    .A1(net147),
    .A2(net245),
    .A3(net14),
    .S0(net998),
    .S1(net758),
    .X(net261));
 sky130_fd_sc_hd__mux4_2 c335 (.A0(net862),
    .A1(net258),
    .A2(net1034),
    .A3(net1004),
    .S0(net1006),
    .S1(net764),
    .X(net262));
 sky130_fd_sc_hd__mux4_1 c336 (.A0(net258),
    .A1(net248),
    .A2(net121),
    .A3(net977),
    .S0(net1023),
    .S1(net758),
    .X(net263));
 sky130_fd_sc_hd__a2111o_1 c337 (.A1(net6),
    .A2(net119),
    .B1(net686),
    .C1(clknet_1_1__leaf_net768),
    .D1(net769),
    .X(net264));
 sky130_fd_sc_hd__mux4_1 c338 (.A0(net132),
    .A1(net141),
    .A2(net258),
    .A3(net130),
    .S0(net1050),
    .S1(net769),
    .X(net265));
 sky130_fd_sc_hd__mux4_1 c339 (.A0(net862),
    .A1(net253),
    .A2(net686),
    .A3(net1008),
    .S0(net726),
    .S1(net949),
    .X(net266));
 sky130_fd_sc_hd__mux4_1 c340 (.A0(net218),
    .A1(net104),
    .A2(net262),
    .A3(net902),
    .S0(net949),
    .S1(clknet_1_1__leaf_net768),
    .X(net267));
 sky130_fd_sc_hd__mux4_1 c341 (.A0(net261),
    .A1(net234),
    .A2(net998),
    .A3(net1050),
    .S0(net1044),
    .S1(net700),
    .X(net268));
 sky130_fd_sc_hd__mux4_1 c342 (.A0(net104),
    .A1(clknet_1_1__leaf_net264),
    .A2(net258),
    .A3(net968),
    .S0(net1026),
    .S1(clknet_1_1__leaf_net768),
    .X(net269));
 sky130_fd_sc_hd__a2111o_1 c343 (.A1(net224),
    .A2(net888),
    .B1(net258),
    .C1(net1104),
    .D1(clknet_1_0__leaf_net264),
    .X(net270));
 sky130_fd_sc_hd__mux4_1 c344 (.A0(clknet_1_1__leaf_net254),
    .A1(net726),
    .A2(net769),
    .A3(net771),
    .S0(net773),
    .S1(net945),
    .X(net271));
 sky130_fd_sc_hd__mux4_1 c345 (.A0(net879),
    .A1(clknet_1_0__leaf_net269),
    .A2(net258),
    .A3(net700),
    .S0(clknet_1_0__leaf_net768),
    .S1(net775),
    .X(net272));
 sky130_fd_sc_hd__mux4_1 c346 (.A0(net262),
    .A1(net993),
    .A2(net258),
    .A3(clknet_1_0__leaf_net768),
    .S0(net774),
    .S1(net945),
    .X(net273));
 sky130_fd_sc_hd__mux4_1 c347 (.A0(net262),
    .A1(net685),
    .A2(net726),
    .A3(net769),
    .S0(net774),
    .S1(net775),
    .X(net274));
 sky130_fd_sc_hd__mux4_1 c348 (.A0(net93),
    .A1(net862),
    .A2(net1037),
    .A3(net1058),
    .S0(clknet_1_0__leaf_net767),
    .S1(net776),
    .X(net275));
 sky130_fd_sc_hd__mux4_1 c349 (.A0(net902),
    .A1(net224),
    .A2(net258),
    .A3(clknet_1_0__leaf_net269),
    .S0(net945),
    .S1(net775),
    .X(net276));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(net137),
    .A1(net121),
    .A2(net710),
    .A3(net712),
    .S0(net775),
    .S1(net776),
    .X(net277));
 sky130_fd_sc_hd__a2111o_1 c351 (.A1(net245),
    .A2(net236),
    .B1(clknet_1_0__leaf_net269),
    .C1(net261),
    .D1(net726),
    .X(net278));
 sky130_fd_sc_hd__mux4_1 c352 (.A0(net870),
    .A1(net46),
    .A2(net236),
    .A3(net81),
    .S0(net967),
    .S1(net685),
    .X(net279));
 sky130_fd_sc_hd__mux4_1 c353 (.A0(net968),
    .A1(net87),
    .A2(clknet_1_0__leaf_net232),
    .A3(net134),
    .S0(net686),
    .S1(net773),
    .X(net280));
 sky130_fd_sc_hd__mux4_1 c354 (.A0(net130),
    .A1(net903),
    .A2(net1029),
    .A3(net972),
    .S0(net968),
    .S1(net685),
    .X(net281));
 sky130_fd_sc_hd__mux4_2 c355 (.A0(net281),
    .A1(net888),
    .A2(net870),
    .A3(net163),
    .S0(net971),
    .S1(net752),
    .X(net282));
 sky130_fd_sc_hd__mux4_2 c356 (.A0(net153),
    .A1(net201),
    .A2(net34),
    .A3(net1029),
    .S0(net1076),
    .S1(net765),
    .X(net283));
 sky130_fd_sc_hd__mux4_2 c357 (.A0(net1055),
    .A1(net34),
    .A2(net1044),
    .A3(net971),
    .S0(net690),
    .S1(net771),
    .X(net284));
 sky130_fd_sc_hd__mux4_2 c358 (.A0(net1104),
    .A1(net1035),
    .A2(net1010),
    .A3(net130),
    .S0(net46),
    .S1(net718),
    .X(net285));
 sky130_fd_sc_hd__mux4_2 c359 (.A0(net134),
    .A1(net879),
    .A2(net283),
    .A3(net1070),
    .S0(net284),
    .S1(net690),
    .X(net955));
 sky130_fd_sc_hd__mux4_1 c360 (.A0(net146),
    .A1(net1104),
    .A2(net1021),
    .A3(net283),
    .S0(net134),
    .S1(net718),
    .X(net286));
 sky130_fd_sc_hd__mux4_1 c361 (.A0(net34),
    .A1(net988),
    .A2(net968),
    .A3(net1033),
    .S0(net279),
    .S1(net1029),
    .X(net287));
 sky130_fd_sc_hd__mux4_2 c362 (.A0(net68),
    .A1(net153),
    .A2(net1089),
    .A3(net281),
    .S0(net752),
    .S1(net765),
    .X(net288));
 sky130_fd_sc_hd__mux4_1 c363 (.A0(net140),
    .A1(net1083),
    .A2(net870),
    .A3(net965),
    .S0(net248),
    .S1(net235),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 c364 (.A0(net1126),
    .A1(clknet_1_0__leaf_net280),
    .A2(net169),
    .A3(net284),
    .S0(net1021),
    .S1(net1005),
    .X(net290));
 sky130_fd_sc_hd__mux4_1 c365 (.A0(net287),
    .A1(clknet_1_0__leaf_net232),
    .A2(net1048),
    .A3(net672),
    .S0(net1006),
    .S1(net1005),
    .X(net291));
 sky130_fd_sc_hd__mux4_1 c366 (.A0(clknet_1_1__leaf_net280),
    .A1(net169),
    .A2(net202),
    .A3(net1069),
    .S0(net1005),
    .S1(net779),
    .X(net292));
 sky130_fd_sc_hd__mux4_1 c367 (.A0(net279),
    .A1(clknet_1_0__leaf_net269),
    .A2(net1126),
    .A3(net1084),
    .S0(net672),
    .S1(net1005),
    .X(net293));
 sky130_fd_sc_hd__mux4_1 c368 (.A0(net1082),
    .A1(net955),
    .A2(net285),
    .A3(net139),
    .S0(net1005),
    .S1(net781),
    .X(net294));
 sky130_fd_sc_hd__mux4_1 c369 (.A0(net282),
    .A1(net294),
    .A2(net1045),
    .A3(net39),
    .S0(net1006),
    .S1(net1005),
    .X(net295));
 sky130_fd_sc_hd__mux4_2 c370 (.A0(net975),
    .A1(net281),
    .A2(net1107),
    .A3(net1071),
    .S0(net956),
    .S1(net945),
    .X(net296));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(net294),
    .A1(net46),
    .A2(net968),
    .A3(net1),
    .S0(net296),
    .S1(net1005),
    .X(net297));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net1072),
    .A1(net294),
    .A2(net1042),
    .A3(clknet_1_1__leaf_net948),
    .S0(net1006),
    .S1(net1005),
    .X(net298));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net968),
    .A1(net155),
    .A2(net1039),
    .A3(clknet_1_1__leaf_net948),
    .S0(net1005),
    .S1(net781),
    .X(net299));
 sky130_fd_sc_hd__mux4_1 c374 (.A0(net253),
    .A1(net181),
    .A2(net1056),
    .A3(net1021),
    .S0(net50),
    .S1(net988),
    .X(net300));
 sky130_fd_sc_hd__mux4_1 c375 (.A0(net287),
    .A1(net857),
    .A2(net942),
    .A3(net61),
    .S0(net1089),
    .S1(net752),
    .X(net301));
 sky130_fd_sc_hd__mux4_1 c376 (.A0(net50),
    .A1(net1053),
    .A2(net1033),
    .A3(net1012),
    .S0(net1020),
    .S1(net783),
    .X(net302));
 sky130_fd_sc_hd__mux4_1 c377 (.A0(net882),
    .A1(net861),
    .A2(net1021),
    .A3(net302),
    .S0(net857),
    .S1(clknet_1_1__leaf_net930),
    .X(net303));
 sky130_fd_sc_hd__mux4_2 c378 (.A0(net1014),
    .A1(net967),
    .A2(net1045),
    .A3(net700),
    .S0(net765),
    .S1(net783),
    .X(net304));
 sky130_fd_sc_hd__mux4_2 c379 (.A0(net285),
    .A1(net50),
    .A2(net861),
    .A3(net1009),
    .S0(net935),
    .S1(net782),
    .X(net305));
 sky130_fd_sc_hd__mux4_1 c380 (.A0(net1056),
    .A1(net1039),
    .A2(net181),
    .A3(net1014),
    .S0(net940),
    .S1(net783),
    .X(net306));
 sky130_fd_sc_hd__mux4_1 c381 (.A0(net861),
    .A1(net306),
    .A2(net304),
    .A3(net1056),
    .S0(net955),
    .S1(net1008),
    .X(net307));
 sky130_fd_sc_hd__mux4_1 c382 (.A0(net234),
    .A1(net181),
    .A2(net55),
    .A3(net1008),
    .S0(net752),
    .S1(clknet_1_1__leaf_net925),
    .X(net953));
 sky130_fd_sc_hd__mux4_1 c383 (.A0(net1045),
    .A1(net0),
    .A2(net882),
    .A3(clknet_1_0__leaf_net953),
    .S0(net1028),
    .S1(net752),
    .X(net308));
 sky130_fd_sc_hd__mux4_1 c384 (.A0(net1033),
    .A1(net201),
    .A2(net1045),
    .A3(net965),
    .S0(net181),
    .S1(clknet_1_1__leaf_net953),
    .X(net309));
 sky130_fd_sc_hd__mux4_1 c385 (.A0(net860),
    .A1(net303),
    .A2(net943),
    .A3(clknet_1_1__leaf_net308),
    .S0(net304),
    .S1(clknet_1_0__leaf_net953),
    .X(net310));
 sky130_fd_sc_hd__mux4_2 c386 (.A0(net305),
    .A1(clknet_1_0__leaf_net308),
    .A2(net908),
    .A3(clknet_1_0__leaf_net953),
    .S0(clknet_1_1__leaf_net930),
    .S1(net988),
    .X(net311));
 sky130_fd_sc_hd__mux4_2 c387 (.A0(clknet_1_0__leaf_net232),
    .A1(net311),
    .A2(net1035),
    .A3(net967),
    .S0(net1012),
    .S1(net940),
    .X(net952));
 sky130_fd_sc_hd__mux4_1 c388 (.A0(net1081),
    .A1(net860),
    .A2(net302),
    .A3(net284),
    .S0(clknet_1_0__leaf_net953),
    .S1(net945),
    .X(net926));
 sky130_fd_sc_hd__mux4_2 c389 (.A0(net284),
    .A1(net135),
    .A2(clknet_1_1__leaf_net952),
    .A3(net1039),
    .S0(net1052),
    .S1(net1021),
    .X(net312));
 sky130_fd_sc_hd__mux4_1 c390 (.A0(net61),
    .A1(net304),
    .A2(net284),
    .A3(net253),
    .S0(net181),
    .S1(clknet_1_1__leaf_net925),
    .X(net313));
 sky130_fd_sc_hd__mux4_1 c391 (.A0(net946),
    .A1(clknet_1_1__leaf_net953),
    .A2(net1081),
    .A3(net698),
    .S0(clknet_1_0__leaf_net948),
    .S1(net935),
    .X(net314));
 sky130_fd_sc_hd__mux4_1 c392 (.A0(clknet_1_1__leaf_net182),
    .A1(net908),
    .A2(clknet_1_0__leaf_net952),
    .A3(clknet_1_1__leaf_net953),
    .S0(net738),
    .S1(net758),
    .X(net315));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net314),
    .A1(net67),
    .A2(net863),
    .A3(net1045),
    .S0(net700),
    .S1(net949),
    .X(net316));
 sky130_fd_sc_hd__mux4_1 c394 (.A0(net302),
    .A1(net170),
    .A2(clknet_1_0__leaf_net316),
    .A3(clknet_1_1__leaf_net953),
    .S0(net698),
    .S1(net949),
    .X(net317));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net136),
    .A1(clknet_1_1__leaf_net316),
    .A2(net988),
    .A3(net967),
    .S0(net751),
    .S1(net758),
    .X(net318));
 sky130_fd_sc_hd__and3_2 c396 (.A(net1042),
    .B(net79),
    .C(net87),
    .X(net319));
 sky130_fd_sc_hd__and3_4 c397 (.A(net1031),
    .B(net74),
    .C(net213),
    .X(net320));
 sky130_fd_sc_hd__and3_4 c398 (.A(net1018),
    .B(net79),
    .C(net992),
    .X(net321));
 sky130_fd_sc_hd__and3_1 c399 (.A(net990),
    .B(net1043),
    .C(net207),
    .X(net322));
 sky130_fd_sc_hd__and2_2 c400 (.A(net195),
    .B(net1091),
    .X(net323));
 sky130_fd_sc_hd__and3_1 c401 (.A(net207),
    .B(net212),
    .C(net1091),
    .X(net324));
 sky130_fd_sc_hd__and3_1 c402 (.A(net68),
    .B(net79),
    .C(net982),
    .X(net325));
 sky130_fd_sc_hd__a2111o_4 c403 (.A1(net982),
    .A2(net322),
    .B1(net211),
    .C1(net1000),
    .D1(net75),
    .X(net326));
 sky130_fd_sc_hd__and3_4 c404 (.A(net608),
    .B(net320),
    .C(net321),
    .X(net327));
 sky130_fd_sc_hd__and3_1 c405 (.A(net211),
    .B(net1000),
    .C(net996),
    .X(net328));
 sky130_fd_sc_hd__a2111o_4 c406 (.A1(net997),
    .A2(net195),
    .B1(net203),
    .C1(net328),
    .D1(net1043),
    .X(net329));
 sky130_fd_sc_hd__and3_1 c407 (.A(net195),
    .B(net211),
    .C(net903),
    .X(net330));
 sky130_fd_sc_hd__a2111o_2 c408 (.A1(net329),
    .A2(net326),
    .B1(net330),
    .C1(net322),
    .D1(net324),
    .X(net331));
 sky130_fd_sc_hd__a2111o_1 c409 (.A1(net321),
    .A2(net331),
    .B1(net324),
    .C1(net327),
    .D1(net82),
    .X(net332));
 sky130_fd_sc_hd__and3_2 c410 (.A(net328),
    .B(net1000),
    .C(net867),
    .X(net333));
 sky130_fd_sc_hd__sdfbbn_2 c411 (.CLK_N(clknet_4_8_0_clk),
    .D(net327),
    .RESET_B(net333),
    .SCD(net982),
    .SCE(net198),
    .SET_B(net657),
    .Q(net335),
    .Q_N(net334));
 sky130_fd_sc_hd__mux4_2 c412 (.A0(net330),
    .A1(net325),
    .A2(net335),
    .A3(net212),
    .S0(net1106),
    .S1(net1017),
    .X(net336));
 sky130_fd_sc_hd__and3_4 c413 (.A(net333),
    .B(net331),
    .C(net321),
    .X(net959));
 sky130_fd_sc_hd__mux4_1 c414 (.A0(net322),
    .A1(net324),
    .A2(net964),
    .A3(net1017),
    .S0(net75),
    .S1(net333),
    .X(net337));
 sky130_fd_sc_hd__dfbbn_2 c415 (.CLK_N(clknet_4_10_0_clk),
    .D(net331),
    .RESET_B(net327),
    .SET_B(net656),
    .Q(net339),
    .Q_N(net338));
 sky130_fd_sc_hd__or4bb_2 c416 (.A(net335),
    .B(net212),
    .C_N(net338),
    .D_N(net657),
    .X(net340));
 sky130_fd_sc_hd__mux4_2 c417 (.A0(net325),
    .A1(net333),
    .A2(net966),
    .A3(net982),
    .S0(net338),
    .S1(net657),
    .X(net341));
 sky130_fd_sc_hd__a2111o_1 c418 (.A1(net77),
    .A2(net329),
    .B1(net979),
    .C1(net657),
    .D1(net1006),
    .X(net342));
 sky130_fd_sc_hd__a2111o_1 c419 (.A1(net333),
    .A2(net103),
    .B1(net96),
    .C1(net200),
    .D1(clknet_1_1__leaf_net230),
    .X(net343));
 sky130_fd_sc_hd__mux4_1 c420 (.A0(net965),
    .A1(net1047),
    .A2(net996),
    .A3(net1044),
    .S0(net979),
    .S1(net1007),
    .X(net344));
 sky130_fd_sc_hd__sdfbbn_2 c421 (.CLK_N(clknet_4_8_0_clk),
    .D(net203),
    .RESET_B(net1098),
    .SCD(net1011),
    .SCE(net1047),
    .SET_B(net964),
    .Q(net346),
    .Q_N(net345));
 sky130_fd_sc_hd__mux4_2 c422 (.A0(net200),
    .A1(net221),
    .A2(net864),
    .A3(net209),
    .S0(net345),
    .S1(net1008),
    .X(net347));
 sky130_fd_sc_hd__mux4_2 c423 (.A0(net196),
    .A1(net333),
    .A2(net325),
    .A3(net1047),
    .S0(net974),
    .S1(net969),
    .X(net348));
 sky130_fd_sc_hd__a2111o_1 c424 (.A1(net220),
    .A2(net1062),
    .B1(clknet_1_0__leaf_net343),
    .C1(net221),
    .D1(net657),
    .X(net349));
 sky130_fd_sc_hd__mux4_1 c425 (.A0(net203),
    .A1(net1083),
    .A2(clknet_1_0__leaf_net343),
    .A3(net965),
    .S0(net876),
    .S1(net979),
    .X(net350));
 sky130_fd_sc_hd__a2111o_1 c426 (.A1(net324),
    .A2(net957),
    .B1(clknet_1_0__leaf_net343),
    .C1(net220),
    .D1(net327),
    .X(net351));
 sky130_fd_sc_hd__a2111o_1 c427 (.A1(net346),
    .A2(clknet_1_0__leaf_net343),
    .B1(net347),
    .C1(net972),
    .D1(net348),
    .X(net352));
 sky130_fd_sc_hd__mux4_2 c428 (.A0(net1122),
    .A1(net1064),
    .A2(net1036),
    .A3(net342),
    .S0(net336),
    .S1(net1092),
    .X(net353));
 sky130_fd_sc_hd__a2111o_1 c429 (.A1(net325),
    .A2(net969),
    .B1(clknet_1_0__leaf_net343),
    .C1(net979),
    .D1(net1063),
    .X(net354));
 sky130_fd_sc_hd__mux4_1 c430 (.A0(net1047),
    .A1(net346),
    .A2(net1083),
    .A3(clknet_1_0__leaf_net343),
    .S0(net221),
    .S1(net327),
    .X(net355));
 sky130_fd_sc_hd__mux4_1 c431 (.A0(net903),
    .A1(clknet_1_1__leaf_net230),
    .A2(net329),
    .A3(clknet_1_0__leaf_net354),
    .S0(clknet_1_1__leaf_net232),
    .S1(net348),
    .X(net356));
 sky130_fd_sc_hd__sdfbbp_1 c432 (.CLK(clknet_4_9_0_clk),
    .D(clknet_1_0__leaf_net354),
    .RESET_B(net215),
    .SCD(net334),
    .SCE(net345),
    .SET_B(net219),
    .Q(net358),
    .Q_N(net357));
 sky130_fd_sc_hd__mux4_1 c433 (.A0(net214),
    .A1(clknet_1_0__leaf_net354),
    .A2(net357),
    .A3(net859),
    .S0(net869),
    .S1(net676),
    .X(net359));
 sky130_fd_sc_hd__mux4_1 c434 (.A0(clknet_1_1__leaf_net232),
    .A1(net982),
    .A2(clknet_1_0__leaf_net354),
    .A3(net996),
    .S0(net864),
    .S1(net1008),
    .X(net360));
 sky130_fd_sc_hd__mux4_1 c435 (.A0(net328),
    .A1(net73),
    .A2(net676),
    .A3(clknet_1_1__leaf_net706),
    .S0(net785),
    .S1(clknet_1_1__leaf_net951),
    .X(net361));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net864),
    .A1(clknet_1_0__leaf_net354),
    .A2(net347),
    .A3(net76),
    .S0(net1067),
    .S1(clknet_1_0__leaf_net951),
    .X(net362));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(clknet_1_0__leaf_net361),
    .A1(net215),
    .A2(net357),
    .A3(clknet_1_0__leaf_net354),
    .S0(net784),
    .S1(clknet_1_0__leaf_net787),
    .X(net363));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(clknet_1_0__leaf_net361),
    .A1(clknet_1_0__leaf_net354),
    .A2(net198),
    .A3(net1090),
    .S0(net329),
    .S1(clknet_1_0__leaf_net951),
    .X(net364));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net358),
    .A1(net209),
    .A2(clknet_1_0__leaf_net706),
    .A3(clknet_1_1__leaf_net767),
    .S0(net788),
    .S1(net790),
    .X(net365));
 sky130_fd_sc_hd__mux4_2 c440 (.A0(clknet_1_1__leaf_net365),
    .A1(net116),
    .A2(net966),
    .A3(net1013),
    .S0(clknet_1_0__leaf_net706),
    .S1(clknet_1_1__leaf_net767),
    .X(net913));
 sky130_fd_sc_hd__a2111o_1 c441 (.A1(net110),
    .A2(clknet_1_0__leaf_net343),
    .B1(net321),
    .C1(net334),
    .D1(net1008),
    .X(net366));
 sky130_fd_sc_hd__a2111o_1 c442 (.A1(net216),
    .A2(net213),
    .B1(net977),
    .C1(net235),
    .D1(net904),
    .X(net367));
 sky130_fd_sc_hd__a2111o_1 c443 (.A1(net1023),
    .A2(net891),
    .B1(net358),
    .C1(net1104),
    .D1(net117),
    .X(net368));
 sky130_fd_sc_hd__sdfbbn_1 c444 (.CLK_N(clknet_4_9_0_clk),
    .D(net367),
    .RESET_B(net116),
    .SCD(net85),
    .SCE(clknet_1_1__leaf_net366),
    .SET_B(net347),
    .Q(net370),
    .Q_N(net369));
 sky130_fd_sc_hd__mux4_1 c445 (.A0(clknet_1_0__leaf_net366),
    .A1(net967),
    .A2(net119),
    .A3(net197),
    .S0(clknet_1_1__leaf_net232),
    .S1(net1020),
    .X(net371));
 sky130_fd_sc_hd__mux4_1 c446 (.A0(net1066),
    .A1(net980),
    .A2(net239),
    .A3(net972),
    .S0(clknet_1_1__leaf_net913),
    .S1(clknet_1_1__leaf_net787),
    .X(net372));
 sky130_fd_sc_hd__a2111o_4 c447 (.A1(net215),
    .A2(net336),
    .B1(net977),
    .C1(net984),
    .D1(net1008),
    .X(net919));
 sky130_fd_sc_hd__mux4_1 c448 (.A0(net116),
    .A1(net886),
    .A2(net369),
    .A3(net1042),
    .S0(net235),
    .S1(net1004),
    .X(net373));
 sky130_fd_sc_hd__a2111o_1 c449 (.A1(net373),
    .A2(net327),
    .B1(clknet_1_0__leaf_net913),
    .C1(net238),
    .D1(net686),
    .X(net374));
 sky130_fd_sc_hd__mux4_1 c450 (.A0(net243),
    .A1(net357),
    .A2(net970),
    .A3(net244),
    .S0(net369),
    .S1(net1008),
    .X(net375));
 sky130_fd_sc_hd__a2111o_1 c451 (.A1(net373),
    .A2(net375),
    .B1(net370),
    .C1(net957),
    .D1(net995),
    .X(net376));
 sky130_fd_sc_hd__mux4_1 c452 (.A0(net964),
    .A1(net238),
    .A2(net116),
    .A3(net980),
    .S0(net666),
    .S1(net1008),
    .X(net377));
 sky130_fd_sc_hd__a2111o_1 c453 (.A1(net335),
    .A2(net68),
    .B1(net246),
    .C1(net1029),
    .D1(clknet_1_1__leaf_net913),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 c454 (.A0(clknet_1_1__leaf_net230),
    .A1(net114),
    .A2(net1011),
    .A3(net368),
    .S0(net931),
    .S1(net693),
    .X(net379));
 sky130_fd_sc_hd__a2111o_1 c455 (.A1(net1030),
    .A2(net975),
    .B1(net666),
    .C1(net734),
    .D1(clknet_1_0__leaf_net787),
    .X(net380));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(net375),
    .A1(net887),
    .A2(net334),
    .A3(net972),
    .S0(net919),
    .S1(net980),
    .X(net381));
 sky130_fd_sc_hd__a2111o_2 c457 (.A1(net243),
    .A2(net367),
    .B1(net975),
    .C1(net866),
    .D1(net682),
    .X(net382));
 sky130_fd_sc_hd__a2111o_1 c458 (.A1(net368),
    .A2(net382),
    .B1(clknet_1_0__leaf_net378),
    .C1(net676),
    .D1(net737),
    .X(net383));
 sky130_fd_sc_hd__mux4_2 c459 (.A0(net209),
    .A1(net977),
    .A2(net320),
    .A3(net335),
    .S0(net848),
    .S1(net357),
    .X(net944));
 sky130_fd_sc_hd__sdfrbp_1 c460 (.CLK(clknet_4_9_0_clk),
    .D(net382),
    .RESET_B(net334),
    .SCD(net984),
    .SCE(net1100),
    .Q(net385),
    .Q_N(net384));
 sky130_fd_sc_hd__a2111o_1 c461 (.A1(net382),
    .A2(net385),
    .B1(net345),
    .C1(net1100),
    .D1(clknet_1_1__leaf_net767),
    .X(net386));
 sky130_fd_sc_hd__mux4_1 c462 (.A0(clknet_1_0__leaf_net233),
    .A1(net1104),
    .A2(net946),
    .A3(net21),
    .S0(net1035),
    .S1(net685),
    .X(net387));
 sky130_fd_sc_hd__mux4_1 c463 (.A0(clknet_1_0__leaf_net372),
    .A1(net1010),
    .A2(net21),
    .A3(net966),
    .S0(clknet_1_1__leaf_net232),
    .S1(net202),
    .X(net388));
 sky130_fd_sc_hd__mux4_1 c464 (.A0(clknet_1_0__leaf_net913),
    .A1(clknet_1_1__leaf_net343),
    .A2(net202),
    .A3(net1107),
    .S0(clknet_1_0__leaf_net767),
    .S1(clknet_1_0__leaf_net768),
    .X(net389));
 sky130_fd_sc_hd__mux4_1 c465 (.A0(net241),
    .A1(net114),
    .A2(net358),
    .A3(clknet_1_1__leaf_net343),
    .S0(net1039),
    .S1(net773),
    .X(net390));
 sky130_fd_sc_hd__mux4_1 c466 (.A0(net390),
    .A1(clknet_1_0__leaf_net275),
    .A2(net1089),
    .A3(net879),
    .S0(net1009),
    .S1(net791),
    .X(net391));
 sky130_fd_sc_hd__mux4_1 c467 (.A0(net1074),
    .A1(clknet_1_1__leaf_net343),
    .A2(net919),
    .A3(clknet_1_0__leaf_net706),
    .S0(net945),
    .S1(net776),
    .X(net392));
 sky130_fd_sc_hd__mux4_2 c468 (.A0(net348),
    .A1(net946),
    .A2(net1010),
    .A3(net1032),
    .S0(net23),
    .S1(net775),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 c469 (.A0(net119),
    .A1(net194),
    .A2(net1039),
    .A3(net1022),
    .S0(clknet_1_1__leaf_net372),
    .S1(net741),
    .X(net394));
 sky130_fd_sc_hd__mux4_1 c470 (.A0(net87),
    .A1(net1016),
    .A2(net879),
    .A3(clknet_1_0__leaf_net269),
    .S0(net709),
    .S1(net775),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 c471 (.A0(net1022),
    .A1(net859),
    .A2(net919),
    .A3(net1084),
    .S0(clknet_1_0__leaf_net767),
    .S1(net775),
    .X(net396));
 sky130_fd_sc_hd__mux4_1 c472 (.A0(clknet_1_0__leaf_net396),
    .A1(net897),
    .A2(clknet_1_1__leaf_net233),
    .A3(net919),
    .S0(clknet_1_0__leaf_net269),
    .S1(net1037),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(net347),
    .A1(net1083),
    .A2(clknet_1_1__leaf_net343),
    .A3(net919),
    .S0(clknet_1_1__leaf_net768),
    .S1(net792),
    .X(net398));
 sky130_fd_sc_hd__mux4_1 c474 (.A0(net995),
    .A1(net984),
    .A2(clknet_1_0__leaf_net380),
    .A3(clknet_1_1__leaf_net913),
    .S0(net690),
    .S1(net941),
    .X(net399));
 sky130_fd_sc_hd__mux4_2 c475 (.A0(net370),
    .A1(net241),
    .A2(net966),
    .A3(clknet_1_0__leaf_net380),
    .S0(net764),
    .S1(net928),
    .X(net400));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(net193),
    .A1(clknet_1_1__leaf_net233),
    .A2(clknet_1_1__leaf_net232),
    .A3(clknet_1_1__leaf_net396),
    .S0(net82),
    .S1(net928),
    .X(net401));
 sky130_fd_sc_hd__mux4_1 c477 (.A0(net966),
    .A1(net320),
    .A2(net193),
    .A3(net1044),
    .S0(net676),
    .S1(net928),
    .X(net402));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(net897),
    .A1(net975),
    .A2(net1034),
    .A3(net857),
    .S0(net793),
    .S1(net928),
    .X(net403));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(net403),
    .A1(net973),
    .A2(clknet_1_0__leaf_net380),
    .A3(net1044),
    .S0(net774),
    .S1(net928),
    .X(net404));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net402),
    .A1(net404),
    .A2(net966),
    .A3(clknet_1_0__leaf_net380),
    .S0(net770),
    .S1(net775),
    .X(net405));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(clknet_1_1__leaf_net392),
    .A1(clknet_1_1__leaf_net343),
    .A2(net973),
    .A3(net1044),
    .S0(net393),
    .S1(net776),
    .X(net406));
 sky130_fd_sc_hd__mux4_2 c482 (.A0(net70),
    .A1(net403),
    .A2(net717),
    .A3(net745),
    .S0(net791),
    .S1(net794),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(clknet_1_0__leaf_net399),
    .A1(net407),
    .A2(clknet_1_0__leaf_net392),
    .A3(net792),
    .S0(net928),
    .S1(net794),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c484 (.A0(clknet_1_1__leaf_net389),
    .A1(net1044),
    .A2(net903),
    .A3(net1000),
    .S0(net741),
    .S1(net956),
    .X(net409));
 sky130_fd_sc_hd__mux4_2 c485 (.A0(net1044),
    .A1(net141),
    .A2(net27),
    .A3(net147),
    .S0(net1029),
    .S1(net771),
    .X(net923));
 sky130_fd_sc_hd__mux4_1 c486 (.A0(net1069),
    .A1(net891),
    .A2(net923),
    .A3(net1029),
    .S0(net262),
    .S1(net718),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 c487 (.A0(net891),
    .A1(net320),
    .A2(net1000),
    .A3(net923),
    .S0(net740),
    .S1(net1102),
    .X(net411));
 sky130_fd_sc_hd__mux4_1 c488 (.A0(net888),
    .A1(net33),
    .A2(net248),
    .A3(net31),
    .S0(net770),
    .S1(net795),
    .X(net412));
 sky130_fd_sc_hd__mux4_1 c489 (.A0(clknet_1_0__leaf_net365),
    .A1(net5),
    .A2(net923),
    .A3(net31),
    .S0(net84),
    .S1(net950),
    .X(net413));
 sky130_fd_sc_hd__mux4_1 c490 (.A0(net169),
    .A1(net172),
    .A2(net7),
    .A3(net139),
    .S0(net776),
    .S1(net780),
    .X(net414));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(clknet_1_1__leaf_net343),
    .A1(net414),
    .A2(net1050),
    .A3(net31),
    .S0(net879),
    .S1(net923),
    .X(net415));
 sky130_fd_sc_hd__mux4_1 c492 (.A0(net147),
    .A1(net107),
    .A2(net1023),
    .A3(net972),
    .S0(net865),
    .S1(net68),
    .X(net416));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(net248),
    .A1(net7),
    .A2(net31),
    .A3(net296),
    .S0(clknet_1_1__leaf_net343),
    .S1(net741),
    .X(net417));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(net1042),
    .A1(net1075),
    .A2(net965),
    .A3(net171),
    .S0(net773),
    .S1(net1005),
    .X(net418));
 sky130_fd_sc_hd__mux4_2 c495 (.A0(net320),
    .A1(net1068),
    .A2(net1004),
    .A3(net935),
    .S0(net751),
    .S1(net795),
    .X(net419));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(net194),
    .A1(net1084),
    .A2(net923),
    .A3(net1023),
    .S0(net139),
    .S1(net769),
    .X(net420));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net1004),
    .A1(net685),
    .A2(net924),
    .A3(net945),
    .S0(net778),
    .S1(net795),
    .X(net421));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(net973),
    .A1(net33),
    .A2(net741),
    .A3(net770),
    .S0(net788),
    .S1(net795),
    .X(net422));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(net31),
    .A1(net921),
    .A2(net866),
    .A3(net944),
    .S0(net419),
    .S1(net740),
    .X(net423));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(clknet_1_0__leaf_net913),
    .A1(net422),
    .A2(net923),
    .A3(net908),
    .S0(net686),
    .S1(net738),
    .X(net424));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(net421),
    .A1(net879),
    .A2(net419),
    .A3(net900),
    .S0(net923),
    .S1(net712),
    .X(net425));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(net416),
    .A1(net1000),
    .A2(net31),
    .A3(net923),
    .S0(net237),
    .S1(net750),
    .X(net426));
 sky130_fd_sc_hd__mux4_2 c503 (.A0(net8),
    .A1(net973),
    .A2(net854),
    .A3(net1035),
    .S0(net924),
    .S1(net796),
    .X(net427));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net68),
    .A1(net419),
    .A2(net8),
    .A3(net903),
    .S0(net745),
    .S1(net778),
    .X(net428));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(net155),
    .A1(net419),
    .A2(net27),
    .A3(net745),
    .S1(net777),
    .X(net429));
 sky130_fd_sc_hd__mux4_1 c526 (.A0(net857),
    .A1(net307),
    .A2(net310),
    .A3(clknet_1_0__leaf_net316),
    .S0(net959),
    .S1(net782),
    .X(net430));
 sky130_fd_sc_hd__mux4_1 c527 (.A0(clknet_1_0__leaf_net389),
    .A1(net988),
    .A2(net318),
    .A3(net923),
    .S0(net750),
    .S1(net758),
    .X(net431));
 sky130_fd_sc_hd__and3_1 c528 (.A(net331),
    .B(net326),
    .C(net656),
    .X(net432));
 sky130_fd_sc_hd__buf_1 c529 (.A(net662),
    .X(net433));
 sky130_fd_sc_hd__and3_1 c530 (.A(net330),
    .B(net433),
    .C(net656),
    .X(net434));
 sky130_fd_sc_hd__and3_1 c531 (.A(net1091),
    .B(net341),
    .C(net992),
    .X(net435));
 sky130_fd_sc_hd__buf_1 c532 (.A(net662),
    .X(net436));
 sky130_fd_sc_hd__and2_2 c533 (.A(net433),
    .B(net341),
    .X(net437));
 sky130_fd_sc_hd__and2_2 c534 (.A(net436),
    .B(net205),
    .X(net438));
 sky130_fd_sc_hd__and3_2 c535 (.A(net1042),
    .B(net990),
    .C(net982),
    .X(net439));
 sky130_fd_sc_hd__and3_2 c536 (.A(net434),
    .B(net77),
    .C(net438),
    .X(net440));
 sky130_fd_sc_hd__mux4_1 c537 (.A0(net74),
    .A1(net439),
    .A2(net438),
    .A3(net964),
    .S0(net434),
    .S1(net341),
    .X(net441));
 sky130_fd_sc_hd__and3_1 c538 (.A(net438),
    .B(net330),
    .C(net205),
    .X(net442));
 sky130_fd_sc_hd__and3_2 c539 (.A(net867),
    .B(net442),
    .C(net192),
    .X(net443));
 sky130_fd_sc_hd__and3_2 c540 (.A(net442),
    .B(net438),
    .C(net205),
    .X(net444));
 sky130_fd_sc_hd__mux4_2 c541 (.A0(net341),
    .A1(net213),
    .A2(net330),
    .A3(net198),
    .S0(net433),
    .S1(net439),
    .X(net445));
 sky130_fd_sc_hd__or4bb_1 c542 (.A(net73),
    .B(net331),
    .C_N(net996),
    .D_N(net434),
    .X(net947));
 sky130_fd_sc_hd__sdfbbn_1 c543 (.CLK_N(clknet_4_10_0_clk),
    .D(net322),
    .RESET_B(net436),
    .SCD(net962),
    .SCE(net330),
    .SET_B(net442),
    .Q(net447),
    .Q_N(net446));
 sky130_fd_sc_hd__clkbuf_4 c544 (.A(net661),
    .X(net448));
 sky130_fd_sc_hd__sdfrtn_1 c545 (.CLK_N(clknet_4_10_0_clk),
    .D(net443),
    .RESET_B(net437),
    .SCD(net962),
    .SCE(net434),
    .Q(net449));
 sky130_fd_sc_hd__mux4_2 c546 (.A0(net436),
    .A1(net449),
    .A2(net444),
    .A3(net966),
    .S0(net608),
    .S1(net691),
    .X(net450));
 sky130_fd_sc_hd__or4bb_1 c547 (.A(net449),
    .B(net331),
    .C_N(net1000),
    .D_N(net448),
    .X(net451));
 sky130_fd_sc_hd__mux4_1 c548 (.A0(net443),
    .A1(net451),
    .A2(net962),
    .A3(net439),
    .S0(net449),
    .S1(net989),
    .X(net452));
 sky130_fd_sc_hd__sdfbbp_1 c549 (.CLK(clknet_4_10_0_clk),
    .D(net451),
    .RESET_B(net448),
    .SCD(net434),
    .SCE(net962),
    .SET_B(net1094),
    .Q(net454),
    .Q_N(net453));
 sky130_fd_sc_hd__or4bb_4 c550 (.A(net342),
    .B(net982),
    .C_N(net219),
    .D_N(net676),
    .X(net455));
 sky130_fd_sc_hd__sdfrtp_4 c551 (.CLK(clknet_4_11_0_clk),
    .D(net847),
    .RESET_B(net353),
    .SCD(net961),
    .SCE(net866),
    .Q(net920));
 sky130_fd_sc_hd__sdfbbn_1 c552 (.CLK_N(clknet_4_11_0_clk),
    .D(net961),
    .RESET_B(net920),
    .SCD(net204),
    .SCE(net976),
    .SET_B(net1018),
    .Q(net457),
    .Q_N(net456));
 sky130_fd_sc_hd__a2111o_1 c553 (.A1(net204),
    .A2(clknet_1_1__leaf_net354),
    .B1(net970),
    .C1(net961),
    .D1(net1092),
    .X(net458));
 sky130_fd_sc_hd__mux4_1 c554 (.A0(net447),
    .A1(net454),
    .A2(net336),
    .A3(net456),
    .S0(net961),
    .S1(net799),
    .X(net459));
 sky130_fd_sc_hd__a2111o_1 c555 (.A1(net608),
    .A2(net456),
    .B1(net961),
    .C1(net869),
    .D1(clknet_1_0__leaf_net786),
    .X(net460));
 sky130_fd_sc_hd__a2111o_2 c556 (.A1(net1017),
    .A2(net342),
    .B1(net869),
    .C1(net970),
    .D1(net677),
    .X(net461));
 sky130_fd_sc_hd__a2111o_1 c557 (.A1(net329),
    .A2(net869),
    .B1(net339),
    .C1(net1020),
    .D1(net1018),
    .X(net462));
 sky130_fd_sc_hd__mux4_2 c558 (.A0(net454),
    .A1(net1031),
    .A2(net198),
    .A3(net1022),
    .S0(net462),
    .S1(net677),
    .X(net463));
 sky130_fd_sc_hd__a2111o_4 c559 (.A1(net198),
    .A2(net1105),
    .B1(net1122),
    .C1(net446),
    .D1(net677),
    .X(net464));
 sky130_fd_sc_hd__mux4_1 c560 (.A0(net462),
    .A1(net461),
    .A2(net847),
    .A3(net463),
    .S0(net353),
    .S1(net798),
    .X(net465));
 sky130_fd_sc_hd__a2111o_4 c561 (.A1(net866),
    .A2(net194),
    .B1(net448),
    .C1(net980),
    .D1(net847),
    .X(net466));
 sky130_fd_sc_hd__sdfbbn_1 c562 (.CLK_N(clknet_4_9_0_clk),
    .D(net432),
    .RESET_B(net876),
    .SCD(net1034),
    .SCE(net800),
    .SET_B(net801),
    .Q(net468),
    .Q_N(net467));
 sky130_fd_sc_hd__sdfrtp_1 c563 (.CLK(clknet_4_11_0_clk),
    .D(net451),
    .RESET_B(net961),
    .SCD(net784),
    .SCE(net800),
    .Q(net469));
 sky130_fd_sc_hd__sdfbbp_1 c564 (.CLK(clknet_4_11_0_clk),
    .D(net202),
    .RESET_B(net447),
    .SCD(net432),
    .SCE(net453),
    .SET_B(net961),
    .Q(net471),
    .Q_N(net470));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net1011),
    .A1(net467),
    .A2(net962),
    .A3(net996),
    .S0(net961),
    .S1(net801),
    .X(net472));
 sky130_fd_sc_hd__a2111o_1 c566 (.A1(net339),
    .A2(net438),
    .B1(net970),
    .C1(net462),
    .D1(net799),
    .X(net473));
 sky130_fd_sc_hd__a2111o_1 c567 (.A1(net462),
    .A2(net875),
    .B1(net464),
    .C1(net473),
    .D1(net466),
    .X(net474));
 sky130_fd_sc_hd__or4bb_2 c568 (.A(net219),
    .B(net468),
    .C_N(net972),
    .D_N(net691),
    .X(net934));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(net471),
    .A1(net329),
    .A2(net221),
    .A3(net469),
    .S0(clknet_1_0__leaf_net349),
    .S1(net691),
    .X(net475));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net87),
    .A1(net357),
    .A2(net934),
    .A3(net1037),
    .S0(net801),
    .S1(clknet_1_0__leaf_net803),
    .X(net476));
 sky130_fd_sc_hd__mux4_1 c571 (.A0(net476),
    .A1(net227),
    .A2(net677),
    .A3(net691),
    .S0(net802),
    .S1(clknet_1_0__leaf_net803),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c572 (.A0(net977),
    .A1(net875),
    .A2(net204),
    .A3(net1000),
    .S0(net677),
    .S1(net737),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c573 (.A0(net1090),
    .A1(net448),
    .A2(net227),
    .A3(net244),
    .S0(clknet_1_1__leaf_net380),
    .S1(net326),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c574 (.A0(net247),
    .A1(net384),
    .A2(net973),
    .A3(net1090),
    .S0(net682),
    .S1(net789),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c575 (.A0(net977),
    .A1(net326),
    .A2(clknet_1_1__leaf_net479),
    .A3(clknet_1_1__leaf_net378),
    .S0(net866),
    .S1(net677),
    .X(net481));
 sky130_fd_sc_hd__mux4_1 c576 (.A0(net867),
    .A1(net82),
    .A2(net1004),
    .A3(clknet_1_1__leaf_net479),
    .S0(net244),
    .S1(net712),
    .X(net482));
 sky130_fd_sc_hd__mux4_1 c577 (.A0(net222),
    .A1(net966),
    .A2(net221),
    .A3(clknet_1_0__leaf_net479),
    .S0(net717),
    .S1(net725),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c578 (.A0(net443),
    .A1(net478),
    .A2(clknet_1_1__leaf_net479),
    .A3(net227),
    .S0(clknet_1_1__leaf_net913),
    .S1(clknet_1_1__leaf_net803),
    .X(net484));
 sky130_fd_sc_hd__mux4_1 c579 (.A0(net440),
    .A1(net221),
    .A2(clknet_1_1__leaf_net361),
    .A3(net743),
    .S0(net800),
    .S1(clknet_1_1__leaf_net805),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c580 (.A0(net353),
    .A1(net222),
    .A2(net444),
    .A3(net384),
    .S0(net466),
    .S1(net934),
    .X(net486));
 sky130_fd_sc_hd__mux4_1 c581 (.A0(net980),
    .A1(net962),
    .A2(net443),
    .A3(net437),
    .S0(net345),
    .S1(net676),
    .X(net487));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(clknet_1_1__leaf_net485),
    .A1(net899),
    .A2(net448),
    .A3(net856),
    .S0(net760),
    .S1(clknet_1_1__leaf_net805),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c583 (.A0(clknet_1_0__leaf_net485),
    .A1(clknet_1_0__leaf_net378),
    .A2(net213),
    .A3(net964),
    .S0(net666),
    .S1(net743),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c584 (.A0(net336),
    .A1(net962),
    .A2(net87),
    .S0(clknet_1_1__leaf_net805),
    .S1(net806),
    .X(net490));
 sky130_fd_sc_hd__mux4_1 c585 (.A0(net990),
    .A1(net1030),
    .A2(net238),
    .A3(net732),
    .S0(net801),
    .S1(net1096),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c586 (.A0(net82),
    .A1(net336),
    .A2(net1030),
    .A3(net319),
    .S0(net323),
    .S1(net790),
    .X(net492));
 sky130_fd_sc_hd__mux4_2 c587 (.A0(net469),
    .A1(net934),
    .A2(net899),
    .A3(net323),
    .S0(net807),
    .S1(net810),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c588 (.A0(net469),
    .A1(clknet_1_1__leaf_net479),
    .A2(net107),
    .A3(net734),
    .S0(clknet_1_0__leaf_net805),
    .S1(net809),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c589 (.A0(net437),
    .A1(net1007),
    .A2(clknet_1_1__leaf_net805),
    .A3(net807),
    .S0(net809),
    .S1(net811),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(net899),
    .A1(net493),
    .A2(clknet_1_1__leaf_net380),
    .A3(net1031),
    .S0(net760),
    .S1(net811),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(net492),
    .A1(net444),
    .A2(clknet_1_0__leaf_net349),
    .A3(net733),
    .S0(clknet_1_0__leaf_net804),
    .S1(net810),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c592 (.A0(net919),
    .A1(net492),
    .A2(net715),
    .A3(net717),
    .S0(clknet_1_1__leaf_net803),
    .S1(net811),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(net463),
    .A1(net437),
    .A2(clknet_1_0__leaf_net498),
    .A3(clknet_1_1__leaf_net479),
    .S0(net962),
    .S1(net715),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c594 (.A0(net340),
    .A1(net82),
    .A2(net407),
    .A3(net920),
    .S0(net980),
    .S1(net993),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c595 (.A0(net21),
    .A1(clknet_1_0__leaf_net399),
    .A2(net262),
    .A3(net876),
    .S0(net407),
    .S1(net114),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c596 (.A0(net463),
    .A1(net966),
    .A2(net1017),
    .A3(net971),
    .S0(net809),
    .S1(net812),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c597 (.A0(net886),
    .A1(net878),
    .A2(net454),
    .A3(net964),
    .S0(net762),
    .S1(net808),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c598 (.A0(net876),
    .A1(net407),
    .A2(net1037),
    .A3(net964),
    .S0(net793),
    .S1(net802),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c599 (.A0(clknet_1_1__leaf_net380),
    .A1(net437),
    .A2(clknet_1_1__leaf_net399),
    .A3(net453),
    .S0(net14),
    .S1(net440),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c600 (.A0(net14),
    .A1(net454),
    .A2(net407),
    .A3(net963),
    .S0(net764),
    .S1(net802),
    .X(net506));
 sky130_fd_sc_hd__mux4_2 c601 (.A0(net478),
    .A1(net886),
    .A2(clknet_1_0__leaf_net400),
    .A3(net1022),
    .S0(net921),
    .S1(net851),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(net899),
    .A1(net921),
    .A2(net1004),
    .A3(net935),
    .S0(net812),
    .S1(net813),
    .X(net508));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(net8),
    .A1(net500),
    .A2(net227),
    .A3(net977),
    .S0(clknet_1_0__leaf_net479),
    .S1(net709),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(net16),
    .A1(clknet_1_0__leaf_net399),
    .A2(clknet_1_0__leaf_net507),
    .A3(net758),
    .S0(net811),
    .S1(net813),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(clknet_1_0__leaf_net399),
    .A1(net974),
    .A2(net16),
    .A3(net971),
    .S0(net813),
    .S1(net958),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net920),
    .A1(net980),
    .A2(net974),
    .A3(net690),
    .S0(net710),
    .S1(net812),
    .X(net512));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(clknet_1_1__leaf_net400),
    .A1(net1034),
    .A2(net14),
    .A3(net876),
    .S0(clknet_1_0__leaf_net746),
    .S1(net794),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net961),
    .A1(clknet_1_1__leaf_net507),
    .A2(clknet_1_1__leaf_net380),
    .A3(net937),
    .S0(clknet_1_1__leaf_net269),
    .S1(net744),
    .X(net514));
 sky130_fd_sc_hd__mux4_1 c609 (.A0(clknet_1_0__leaf_net507),
    .A1(net440),
    .A2(net869),
    .A3(net975),
    .S0(net753),
    .S1(net813),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c610 (.A0(clknet_1_1__leaf_net275),
    .A1(net971),
    .A2(net407),
    .A3(net1012),
    .S0(clknet_1_0__leaf_net479),
    .S1(net814),
    .X(net516));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net407),
    .A1(net500),
    .A2(net919),
    .A3(net319),
    .S0(net813),
    .S1(net814),
    .X(net517));
 sky130_fd_sc_hd__mux4_2 c612 (.A0(net974),
    .A1(net358),
    .A2(net723),
    .A3(net812),
    .S0(net958),
    .S1(net814),
    .X(net518));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(clknet_1_1__leaf_net361),
    .A1(net918),
    .A2(net517),
    .A3(clknet_1_0__leaf_net747),
    .S0(net928),
    .S1(net814),
    .X(net519));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(net517),
    .A1(net961),
    .A2(net518),
    .A3(net802),
    .S0(net814),
    .S1(net815),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net512),
    .A1(clknet_1_0__leaf_net507),
    .A2(net966),
    .A3(net744),
    .S0(net753),
    .S1(net814),
    .X(net521));
 sky130_fd_sc_hd__mux4_1 c616 (.A0(net282),
    .A1(net1050),
    .A2(net963),
    .A3(net917),
    .S0(net909),
    .S1(net776),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(net288),
    .A1(net16),
    .A2(net927),
    .A3(net27),
    .S0(net39),
    .S1(net793),
    .X(net523));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(net33),
    .A1(net237),
    .A2(net202),
    .A3(net419),
    .S0(net982),
    .S1(net39),
    .X(net524));
 sky130_fd_sc_hd__mux4_1 c619 (.A0(net82),
    .A1(net106),
    .A2(clknet_1_0__leaf_net299),
    .A3(net283),
    .S0(net963),
    .S1(net771),
    .X(net525));
 sky130_fd_sc_hd__mux4_2 c62 (.A0(net871),
    .A1(net883),
    .A2(net896),
    .A3(net888),
    .S0(net894),
    .S1(net884),
    .X(net0));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net875),
    .A1(net918),
    .A2(net772),
    .A3(net777),
    .S0(net958),
    .S1(net819),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(net321),
    .A1(clknet_1_0__leaf_net913),
    .A2(net296),
    .A3(net1020),
    .S0(net723),
    .S1(net778),
    .X(net527));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(net931),
    .A1(net866),
    .A2(net16),
    .A3(net283),
    .S0(net770),
    .S1(net780),
    .X(net528));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(net973),
    .A1(net18),
    .A2(net427),
    .A3(net119),
    .S0(net467),
    .S1(net754),
    .X(net529));
 sky130_fd_sc_hd__mux4_1 c624 (.A0(net107),
    .A1(net8),
    .A2(net33),
    .A3(net119),
    .S0(net754),
    .S1(net928),
    .X(net530));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net529),
    .A1(net528),
    .A2(net1012),
    .A3(net1031),
    .S0(net1049),
    .S1(net119),
    .X(net531));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net513),
    .A1(net866),
    .A2(net27),
    .A3(net1042),
    .S0(net954),
    .S1(net770),
    .X(net532));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(clknet_1_1__leaf_net299),
    .A1(net296),
    .A2(net107),
    .A3(net762),
    .S0(clknet_1_0__leaf_net805),
    .S1(net922),
    .X(net533));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net468),
    .A1(net1030),
    .A2(net918),
    .A3(net33),
    .S0(net795),
    .S1(clknet_1_0__leaf_net805),
    .X(net534));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(net27),
    .A1(net202),
    .A2(net1000),
    .A3(net33),
    .S0(net763),
    .S1(net938),
    .X(net535));
 sky130_fd_sc_hd__mux4_2 c63 (.A0(net898),
    .A1(net899),
    .A2(net3),
    .A3(net897),
    .S0(net0),
    .S1(net890),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net526),
    .A1(net119),
    .A2(net419),
    .A3(net535),
    .S0(net770),
    .S1(net777),
    .X(net536));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net535),
    .A1(net855),
    .A2(net915),
    .A3(net759),
    .S0(net820),
    .S1(clknet_1_1__leaf_net822),
    .X(net537));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net493),
    .A1(net893),
    .A2(net927),
    .A3(net712),
    .S0(net924),
    .S1(net1101),
    .X(net538));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(clknet_1_0__leaf_net479),
    .A1(net887),
    .A2(net422),
    .A3(clknet_1_0__leaf_net537),
    .S0(net282),
    .S1(net819),
    .X(net539));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net531),
    .A1(net194),
    .A2(net288),
    .A3(net107),
    .S0(net793),
    .S1(clknet_1_0__leaf_net821),
    .X(net540));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net908),
    .A1(net933),
    .A2(net1019),
    .A3(net919),
    .S0(net722),
    .S1(net797),
    .X(net541));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net530),
    .A1(net8),
    .A2(net1030),
    .A3(net725),
    .S0(net772),
    .S1(clknet_1_0__leaf_net821),
    .X(net542));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net541),
    .A1(clknet_1_0__leaf_net542),
    .A2(net933),
    .A3(net954),
    .S0(net759),
    .S1(net817),
    .X(net543));
 sky130_fd_sc_hd__mux4_2 c64 (.A0(net883),
    .A1(net1),
    .A2(net898),
    .A3(net890),
    .S0(net884),
    .S1(net896),
    .X(net2));
 sky130_fd_sc_hd__mux4_2 c65 (.A0(net1027),
    .A1(net871),
    .A2(net881),
    .A3(net880),
    .S0(net1041),
    .S1(net1031),
    .X(net3));
 sky130_fd_sc_hd__and3_2 c66 (.A(net901),
    .B(net1040),
    .C(net890),
    .X(net4));
 sky130_fd_sc_hd__a2111o_1 c660 (.A1(net196),
    .A2(net1036),
    .B1(net86),
    .C1(net75),
    .D1(net691),
    .X(net544));
 sky130_fd_sc_hd__sdfrtp_1 c661 (.CLK(clknet_4_10_0_clk),
    .D(net339),
    .RESET_B(net976),
    .SCD(net858),
    .SCE(net450),
    .Q(net545));
 sky130_fd_sc_hd__a2111o_1 c662 (.A1(net212),
    .A2(net448),
    .B1(net544),
    .C1(net858),
    .D1(net989),
    .X(net546));
 sky130_fd_sc_hd__dlymetal6s2s_1 c663 (.A(net845),
    .X(net547));
 sky130_fd_sc_hd__and3_1 c664 (.A(net79),
    .B(net858),
    .C(net992),
    .X(net548));
 sky130_fd_sc_hd__buf_1 c665 (.A(net844),
    .X(net549));
 sky130_fd_sc_hd__and3_4 c666 (.A(net192),
    .B(net1022),
    .C(net999),
    .X(net911));
 sky130_fd_sc_hd__a2111o_1 c667 (.A1(net548),
    .A2(net546),
    .B1(net544),
    .C1(net999),
    .D1(net547),
    .X(net550));
 sky130_fd_sc_hd__and3_1 c668 (.A(net1036),
    .B(net550),
    .C(net911),
    .X(net551));
 sky130_fd_sc_hd__and3_2 c669 (.A(net69),
    .B(net547),
    .C(net999),
    .X(net552));
 sky130_fd_sc_hd__and3_4 c67 (.A(net1037),
    .B(net879),
    .C(net1025),
    .X(net5));
 sky130_fd_sc_hd__and3_2 c670 (.A(net75),
    .B(net545),
    .C(net453),
    .X(net553));
 sky130_fd_sc_hd__mux4_1 c671 (.A0(net454),
    .A1(net552),
    .A2(net553),
    .A3(net999),
    .S0(net911),
    .S1(net546),
    .X(net554));
 sky130_fd_sc_hd__a2111o_2 c672 (.A1(net1099),
    .A2(net911),
    .B1(net547),
    .C1(net554),
    .D1(net976),
    .X(net555));
 sky130_fd_sc_hd__a2111o_1 c673 (.A1(net858),
    .A2(net552),
    .B1(net1022),
    .C1(net992),
    .D1(net1003),
    .X(net556));
 sky130_fd_sc_hd__buf_2 c674 (.A(net661),
    .X(net557));
 sky130_fd_sc_hd__a2111o_1 c675 (.A1(net205),
    .A2(net545),
    .B1(net444),
    .C1(net553),
    .D1(net999),
    .X(net558));
 sky130_fd_sc_hd__a2111o_1 c676 (.A1(net75),
    .A2(net321),
    .B1(net1097),
    .C1(net445),
    .D1(net999),
    .X(net559));
 sky130_fd_sc_hd__a2111o_1 c677 (.A1(net556),
    .A2(net552),
    .B1(net858),
    .C1(net557),
    .D1(net691),
    .X(net560));
 sky130_fd_sc_hd__a2111o_1 c678 (.A1(net1039),
    .A2(net858),
    .B1(net557),
    .C1(net553),
    .D1(net1003),
    .X(net561));
 sky130_fd_sc_hd__mux4_1 c679 (.A0(net544),
    .A1(net552),
    .A2(net548),
    .A3(net551),
    .S0(net197),
    .S1(net553),
    .X(net562));
 sky130_fd_sc_hd__and3_2 c68 (.A(net1017),
    .B(net883),
    .C(net881),
    .X(net6));
 sky130_fd_sc_hd__a2111o_1 c680 (.A1(net561),
    .A2(net551),
    .B1(net560),
    .C1(net1099),
    .D1(net557),
    .X(net563));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(net553),
    .A1(net556),
    .A2(net435),
    .A3(net561),
    .S0(net548),
    .S1(net665),
    .X(net564));
 sky130_fd_sc_hd__mux4_1 c682 (.A0(net77),
    .A1(net450),
    .A2(net1105),
    .A3(net357),
    .S0(net1016),
    .S1(clknet_1_1__leaf_net706),
    .X(net565));
 sky130_fd_sc_hd__mux4_1 c683 (.A0(net438),
    .A1(net552),
    .A2(net466),
    .A3(net450),
    .S0(net557),
    .S1(net1020),
    .X(net566));
 sky130_fd_sc_hd__mux4_1 c684 (.A0(net554),
    .A1(net1016),
    .A2(net196),
    .A3(clknet_1_0__leaf_net786),
    .S0(net826),
    .S1(net828),
    .X(net567));
 sky130_fd_sc_hd__mux4_1 c685 (.A0(net1108),
    .A1(net444),
    .A2(net552),
    .A3(net557),
    .S0(clknet_1_0__leaf_net477),
    .S1(net1105),
    .X(net568));
 sky130_fd_sc_hd__mux4_1 c686 (.A0(net550),
    .A1(net992),
    .A2(net1105),
    .A3(net1015),
    .S0(clknet_1_1__leaf_net786),
    .S1(net828),
    .X(net569));
 sky130_fd_sc_hd__mux4_1 c687 (.A0(net547),
    .A1(net326),
    .A2(net321),
    .A3(net213),
    .S0(clknet_1_1__leaf_net706),
    .S1(net829),
    .X(net570));
 sky130_fd_sc_hd__mux4_2 c688 (.A0(net69),
    .A1(net550),
    .A2(net326),
    .A3(net1105),
    .S0(net665),
    .S1(net800),
    .X(net571));
 sky130_fd_sc_hd__mux4_1 c689 (.A0(clknet_1_0__leaf_net570),
    .A1(net999),
    .A2(clknet_1_1__leaf_net354),
    .A3(net439),
    .S0(clknet_1_1__leaf_net786),
    .S1(net800),
    .X(net572));
 sky130_fd_sc_hd__a2111o_4 c69 (.A1(net874),
    .A2(net877),
    .B1(net891),
    .C1(net894),
    .D1(net1107),
    .X(net7));
 sky130_fd_sc_hd__mux4_1 c690 (.A0(net551),
    .A1(net339),
    .A2(net553),
    .A3(net221),
    .S0(net85),
    .S1(net824),
    .X(net573));
 sky130_fd_sc_hd__mux4_1 c691 (.A0(net473),
    .A1(net461),
    .A2(net549),
    .A3(net453),
    .S0(net1000),
    .S1(net829),
    .X(net574));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(clknet_1_0__leaf_net477),
    .A1(net560),
    .A2(net86),
    .A3(net338),
    .S0(net557),
    .S1(net828),
    .X(net575));
 sky130_fd_sc_hd__mux4_1 c693 (.A0(clknet_1_1__leaf_net567),
    .A1(net438),
    .A2(clknet_1_0__leaf_net575),
    .A3(net999),
    .S0(net439),
    .S1(net347),
    .X(net576));
 sky130_fd_sc_hd__mux4_1 c694 (.A0(net450),
    .A1(clknet_1_1__leaf_net570),
    .A2(net473),
    .A3(net320),
    .S0(net982),
    .S1(net1039),
    .X(net577));
 sky130_fd_sc_hd__mux4_1 c695 (.A0(net560),
    .A1(net571),
    .A2(net439),
    .A3(net197),
    .S0(net1036),
    .S1(net694),
    .X(net578));
 sky130_fd_sc_hd__mux4_2 c696 (.A0(net558),
    .A1(net1036),
    .A2(net996),
    .A3(net982),
    .S0(net830),
    .S1(net912),
    .X(net579));
 sky130_fd_sc_hd__mux4_1 c697 (.A0(net557),
    .A1(clknet_1_0__leaf_net567),
    .A2(clknet_1_0__leaf_net575),
    .A3(net1036),
    .S0(net552),
    .S1(net830),
    .X(net580));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(net553),
    .A1(clknet_1_1__leaf_net477),
    .A2(net336),
    .A3(net665),
    .S0(net785),
    .S1(net832),
    .X(net581));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(net571),
    .A1(net473),
    .A2(net558),
    .A3(net694),
    .S0(net739),
    .S1(net832),
    .X(net582));
 sky130_fd_sc_hd__or4bb_4 c70 (.A(net1023),
    .B(net874),
    .C_N(net1025),
    .D_N(net6),
    .X(net8));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net554),
    .A1(clknet_1_0__leaf_net570),
    .A2(net555),
    .A3(clknet_1_0__leaf_net581),
    .S0(net799),
    .S1(net832),
    .X(net583));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(net545),
    .A1(net1016),
    .A2(net339),
    .A3(net197),
    .S0(clknet_1_1__leaf_net786),
    .S1(net833),
    .X(net584));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net439),
    .A1(net443),
    .A2(clknet_1_1__leaf_net570),
    .A3(clknet_1_1__leaf_net354),
    .S0(net830),
    .S1(net831),
    .X(net585));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(net547),
    .A1(clknet_1_0__leaf_net581),
    .A2(net739),
    .A3(net755),
    .S0(net830),
    .S1(net831),
    .X(net586));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net385),
    .A1(net1037),
    .A2(net1105),
    .A3(net1036),
    .S0(net887),
    .S1(net1007),
    .X(net587));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(net382),
    .A1(net985),
    .A2(net555),
    .A3(net1019),
    .S0(net753),
    .S1(net831),
    .X(net588));
 sky130_fd_sc_hd__mux4_2 c706 (.A0(net457),
    .A1(net346),
    .A2(net555),
    .A3(net1030),
    .S0(net1095),
    .S1(net830),
    .X(net589));
 sky130_fd_sc_hd__mux4_1 c707 (.A0(net238),
    .A1(net552),
    .A2(net1105),
    .A3(net464),
    .S0(net678),
    .S1(net830),
    .X(net590));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(net443),
    .A1(net382),
    .A2(net455),
    .A3(net964),
    .S0(net832),
    .S1(net837),
    .X(net591));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(net1015),
    .A1(net571),
    .A2(net444),
    .A3(net678),
    .S0(net749),
    .S1(net800),
    .X(net592));
 sky130_fd_sc_hd__and3_1 c71 (.A(net1043),
    .B(net876),
    .C(net879),
    .X(net9));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net326),
    .A1(net584),
    .A2(clknet_1_0__leaf_net568),
    .A3(net1007),
    .S0(net785),
    .S1(net834),
    .X(net593));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net444),
    .A1(clknet_1_1__leaf_net354),
    .A2(clknet_1_0__leaf_net496),
    .A3(net117),
    .S0(net999),
    .S1(net715),
    .X(net594));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(clknet_1_1__leaf_net378),
    .A1(net346),
    .A2(net830),
    .A3(net831),
    .S0(net832),
    .S1(net838),
    .X(net595));
 sky130_fd_sc_hd__mux4_1 c713 (.A0(net552),
    .A1(clknet_1_1__leaf_net581),
    .A2(net440),
    .A3(net466),
    .S0(net1031),
    .S1(net834),
    .X(net596));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(net347),
    .A1(net440),
    .A2(net1036),
    .A3(net964),
    .S0(net694),
    .S1(net907),
    .X(net597));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net546),
    .A1(net893),
    .A2(net466),
    .A3(net1105),
    .S0(net859),
    .S1(net755),
    .X(net598));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net457),
    .A1(net555),
    .A2(net1031),
    .A3(net682),
    .S0(clknet_1_0__leaf_net742),
    .S1(net912),
    .X(net599));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net571),
    .A1(net385),
    .A2(net587),
    .A3(clknet_1_1__leaf_net354),
    .S0(net715),
    .S1(net800),
    .X(net600));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(net244),
    .A1(net213),
    .A2(net464),
    .A3(net682),
    .S0(net749),
    .S1(net829),
    .X(net601));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net964),
    .A1(net470),
    .A2(net846),
    .A3(net689),
    .S0(net839),
    .S1(net840),
    .X(net602));
 sky130_fd_sc_hd__and3_2 c72 (.A(net1024),
    .B(net6),
    .C(net1028),
    .X(net10));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net1022),
    .A1(clknet_1_1__leaf_net498),
    .A2(net1016),
    .A3(net785),
    .S0(net831),
    .S1(clknet_1_0__leaf_net841),
    .X(net603));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net336),
    .A1(net221),
    .A2(net694),
    .A3(net836),
    .S0(net840),
    .S1(clknet_1_1__leaf_net841),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net82),
    .A1(clknet_1_1__leaf_net604),
    .A2(clknet_1_1__leaf_net378),
    .A3(net809),
    .S0(net840),
    .S1(clknet_1_0__leaf_net841),
    .X(net605));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net598),
    .A1(net852),
    .A2(net756),
    .A3(net800),
    .S0(net839),
    .S1(clknet_1_1__leaf_net841),
    .X(net606));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net606),
    .A1(clknet_1_1__leaf_net604),
    .A2(net986),
    .A3(clknet_1_1__leaf_net575),
    .S0(net1007),
    .S1(net840),
    .X(net607));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net246),
    .A1(net327),
    .A2(clknet_1_1__leaf_net604),
    .S0(net756),
    .S1(net840),
    .X(net742));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net859),
    .A1(net1121),
    .A2(net1004),
    .A3(net678),
    .S0(net825),
    .S1(net835),
    .X(net609));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net448),
    .A1(net859),
    .A2(net518),
    .A3(net986),
    .S0(net724),
    .S1(net838),
    .X(net610));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net85),
    .A1(clknet_1_1__leaf_net575),
    .A2(net347),
    .A3(net863),
    .S0(net724),
    .S1(net915),
    .X(net611));
 sky130_fd_sc_hd__mux4_2 c729 (.A0(net464),
    .A1(net117),
    .A2(net244),
    .A3(net986),
    .S0(net1020),
    .S1(net816),
    .X(net612));
 sky130_fd_sc_hd__and3_1 c73 (.A(net881),
    .B(net902),
    .C(net7),
    .X(net11));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net587),
    .A1(net863),
    .A2(net1019),
    .A3(net776),
    .S0(net833),
    .S1(net838),
    .X(net613));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net609),
    .A1(net1121),
    .A2(net358),
    .A3(net612),
    .S0(net688),
    .S1(clknet_1_0__leaf_net742),
    .X(net614));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(net471),
    .A1(net976),
    .A2(net213),
    .A3(net760),
    .S0(net909),
    .S1(net829),
    .X(net615));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(clknet_1_1__leaf_net349),
    .A1(net869),
    .A2(net613),
    .A3(net244),
    .S0(net868),
    .S1(net813),
    .X(net616));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(net393),
    .A1(net117),
    .A2(net262),
    .A3(net464),
    .S0(net772),
    .S1(net813),
    .X(net617));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net213),
    .A1(net615),
    .A2(net986),
    .A3(clknet_1_1__leaf_net913),
    .S0(clknet_1_1__leaf_net804),
    .S1(net834),
    .X(net618));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(net358),
    .A1(net508),
    .A2(net1121),
    .A3(net986),
    .S0(clknet_1_1__leaf_net913),
    .S1(net816),
    .X(net619));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net440),
    .A1(net461),
    .A2(net464),
    .A3(net23),
    .S0(net971),
    .S1(net754),
    .X(net620));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net244),
    .A1(net986),
    .A2(clknet_1_1__leaf_net507),
    .A3(net852),
    .S0(net448),
    .S1(net87),
    .X(net621));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(net601),
    .A1(net321),
    .A2(net868),
    .A3(net745),
    .S0(net909),
    .S1(net825),
    .X(net622));
 sky130_fd_sc_hd__and3_4 c74 (.A(net2),
    .B(net1107),
    .C(net1025),
    .X(net12));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(net518),
    .A1(net587),
    .A2(clknet_1_1__leaf_net349),
    .A3(net470),
    .S0(clknet_1_1__leaf_net569),
    .S1(net683),
    .X(net623));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(net613),
    .A1(net976),
    .A2(net869),
    .A3(net440),
    .S0(clknet_1_1__leaf_net618),
    .S1(net729),
    .X(net624));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(net461),
    .A1(clknet_1_1__leaf_net507),
    .A2(clknet_1_0__leaf_net618),
    .A3(net601),
    .S0(net776),
    .S1(net829),
    .X(net625));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(clknet_1_1__leaf_net568),
    .A1(net963),
    .A2(net393),
    .A3(net794),
    .S0(net958),
    .S1(clknet_1_0__leaf_net843),
    .X(net626));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(clknet_1_1__leaf_net349),
    .A1(clknet_1_1__leaf_net913),
    .A2(net262),
    .A3(net830),
    .S0(clknet_1_0__leaf_net842),
    .S1(clknet_1_0__leaf_net843),
    .X(net627));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(net869),
    .A1(net1022),
    .A2(net612),
    .A3(net859),
    .S0(net739),
    .S1(clknet_1_1__leaf_net842),
    .X(net628));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net555),
    .A1(net619),
    .A2(net849),
    .A3(net960),
    .S0(net835),
    .S1(clknet_1_1__leaf_net843),
    .X(net629));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(net868),
    .A1(net754),
    .A2(net760),
    .A3(net794),
    .S0(net832),
    .S1(clknet_1_0__leaf_net842),
    .X(net630));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net885),
    .A1(net197),
    .A2(net759),
    .A3(net774),
    .S0(clknet_1_0__leaf_net804),
    .S1(net810),
    .X(net631));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net466),
    .A1(net197),
    .A2(net911),
    .A3(clknet_1_1__leaf_net534),
    .S0(clknet_1_1__leaf_net823),
    .S1(net832),
    .X(net632));
 sky130_fd_sc_hd__and2_4 c75 (.A(net12),
    .B(net902),
    .X(net13));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(net859),
    .A1(net1031),
    .A2(net632),
    .A3(net959),
    .S0(clknet_1_1__leaf_net916),
    .S1(clknet_1_1__leaf_net747),
    .X(net633));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net612),
    .A1(net262),
    .A2(clknet_1_1__leaf_net269),
    .A3(net971),
    .S0(net748),
    .S1(clknet_1_1__leaf_net821),
    .X(net634));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(clknet_1_1__leaf_net269),
    .A1(clknet_1_1__leaf_net537),
    .A2(net1019),
    .A3(net1020),
    .S0(clknet_1_1__leaf_net747),
    .S1(net835),
    .X(net635));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(clknet_1_0__leaf_net604),
    .A1(net319),
    .A2(net327),
    .A3(clknet_1_0__leaf_net537),
    .S0(net958),
    .S1(clknet_1_0__leaf_net822),
    .X(net636));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net887),
    .A1(net240),
    .A2(net630),
    .A3(net1039),
    .S0(clknet_1_1__leaf_net269),
    .S1(net776),
    .X(net637));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net999),
    .A1(net631),
    .A2(net39),
    .A3(net717),
    .S0(net753),
    .S1(net795),
    .X(net638));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net114),
    .A1(net1020),
    .A2(net993),
    .A3(net1031),
    .S0(net39),
    .S1(net811),
    .X(net639));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net321),
    .A1(net1058),
    .A2(net893),
    .A3(net772),
    .S0(net818),
    .S1(clknet_1_0__leaf_net823),
    .X(net906));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net1019),
    .A1(net639),
    .A2(net239),
    .A3(net722),
    .S0(net759),
    .S1(net810),
    .X(net640));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net990),
    .A1(net852),
    .A2(clknet_1_0__leaf_net618),
    .A3(net640),
    .S0(net114),
    .S1(net684),
    .X(net641));
 sky130_fd_sc_hd__and2_4 c76 (.A(net880),
    .B(net7),
    .X(net14));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(clknet_1_0__leaf_net569),
    .A1(net610),
    .A2(net39),
    .A3(net852),
    .S0(net757),
    .S1(net827),
    .X(net642));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net172),
    .A1(clknet_1_0__leaf_net498),
    .A2(net905),
    .A3(net638),
    .S0(net327),
    .S1(clknet_1_0__leaf_net916),
    .X(net643));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net893),
    .A1(net1015),
    .A2(net1019),
    .A3(clknet_1_1__leaf_net746),
    .S0(net757),
    .S1(net839),
    .X(net644));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(net323),
    .A1(net1004),
    .A2(net455),
    .A3(net240),
    .S0(net989),
    .X(net707));
 sky130_fd_sc_hd__mux4_1 c764 (.A0(net283),
    .A1(net644),
    .A2(clknet_1_0__leaf_net604),
    .A3(net319),
    .S0(clknet_1_0__leaf_net916),
    .S1(net833),
    .X(net646));
 sky130_fd_sc_hd__mux4_1 c765 (.A0(clknet_1_1__leaf_net496),
    .A1(net733),
    .A2(net740),
    .A3(clknet_1_1__leaf_net746),
    .S0(net763),
    .S1(net827),
    .X(net647));
 sky130_fd_sc_hd__mux4_1 c766 (.A0(net87),
    .A1(net323),
    .A2(net240),
    .A3(net728),
    .S0(clknet_1_1__leaf_net742),
    .S1(net763),
    .X(net648));
 sky130_fd_sc_hd__mux4_1 c767 (.A0(net645),
    .A1(net905),
    .A2(clknet_1_1__leaf_net542),
    .A3(net647),
    .S0(net648),
    .S1(net748),
    .X(net649));
 sky130_fd_sc_hd__mux4_1 c768 (.A0(net1030),
    .A1(net889),
    .A2(net707),
    .A3(net915),
    .S0(net954),
    .S1(net958),
    .X(net650));
 sky130_fd_sc_hd__mux4_1 c769 (.A0(net427),
    .A1(clknet_1_0__leaf_net534),
    .A2(net650),
    .A3(clknet_1_1__leaf_net269),
    .S0(clknet_1_0__leaf_net746),
    .S1(clknet_1_0__leaf_net747),
    .X(net651));
 sky130_fd_sc_hd__and2_2 c77 (.A(net863),
    .B(net1017),
    .X(net15));
 sky130_fd_sc_hd__and2_4 c78 (.A(net15),
    .B(net10),
    .X(net16));
 sky130_fd_sc_hd__a2111o_4 c79 (.A1(net12),
    .A2(net16),
    .B1(net7),
    .C1(net9),
    .D1(net8),
    .X(net17));
 sky130_fd_sc_hd__or4bb_4 c80 (.A(net7),
    .B(net4),
    .C_N(net2),
    .D_N(net15),
    .X(net18));
 sky130_fd_sc_hd__a2111o_4 c81 (.A1(net17),
    .A2(net11),
    .B1(net10),
    .C1(net1042),
    .D1(net1107),
    .X(net19));
 sky130_fd_sc_hd__mux4_2 c82 (.A0(net13),
    .A1(net9),
    .A2(net18),
    .A3(net12),
    .S0(net1016),
    .S1(net11),
    .X(net20));
 sky130_fd_sc_hd__a2111o_4 c83 (.A1(net1034),
    .A2(net15),
    .B1(net1107),
    .C1(net16),
    .D1(net991),
    .X(net21));
 sky130_fd_sc_hd__a2111o_4 c84 (.A1(net9),
    .A2(net17),
    .B1(net1025),
    .C1(net991),
    .D1(net19),
    .X(net22));
 sky130_fd_sc_hd__mux4_2 c85 (.A0(net11),
    .A1(net21),
    .A2(net19),
    .A3(net22),
    .S0(net14),
    .S1(net12),
    .X(net23));
 sky130_fd_sc_hd__a2111o_1 c86 (.A1(net23),
    .A2(net18),
    .B1(net22),
    .C1(net19),
    .D1(net991),
    .X(net24));
 sky130_fd_sc_hd__mux4_2 c87 (.A0(net991),
    .A1(net18),
    .A2(net1107),
    .A3(net23),
    .S0(net887),
    .S1(net987),
    .X(net25));
 sky130_fd_sc_hd__and3_1 c88 (.A(net877),
    .B(net15),
    .C(net1023),
    .X(net26));
 sky130_fd_sc_hd__and3_4 c89 (.A(net1021),
    .B(net882),
    .C(net1024),
    .X(net27));
 sky130_fd_sc_hd__and3_1 c90 (.A(net1),
    .B(net19),
    .C(net1043),
    .X(net28));
 sky130_fd_sc_hd__or4bb_2 c91 (.A(net894),
    .B(net860),
    .C_N(net17),
    .D_N(net1043),
    .X(net29));
 sky130_fd_sc_hd__and3_2 c92 (.A(net4),
    .B(net12),
    .C(net13),
    .X(net30));
 sky130_fd_sc_hd__and3_4 c93 (.A(net28),
    .B(net870),
    .C(net1025),
    .X(net31));
 sky130_fd_sc_hd__a2111o_4 c94 (.A1(net13),
    .A2(net987),
    .B1(net17),
    .C1(net16),
    .D1(net25),
    .X(net32));
 sky130_fd_sc_hd__mux4_2 c95 (.A0(net1023),
    .A1(net874),
    .A2(net28),
    .A3(net1032),
    .S0(net2),
    .S1(net8),
    .X(net33));
 sky130_fd_sc_hd__and3_2 c96 (.A(net890),
    .B(net13),
    .C(net26),
    .X(net34));
 sky130_fd_sc_hd__and3_1 c97 (.A(net17),
    .B(net981),
    .C(net29),
    .X(net35));
 sky130_fd_sc_hd__mux4_2 c98 (.A0(net1018),
    .A1(net35),
    .A2(net981),
    .A3(net4),
    .S0(net27),
    .S1(net28),
    .X(net36));
 sky130_fd_sc_hd__or4bb_4 c99 (.A(net1107),
    .B(net31),
    .C_N(net30),
    .D_N(net981),
    .X(net37));
 sky130_fd_sc_hd__mux4_1 merge790 (.A0(net204),
    .A1(net432),
    .A2(net1003),
    .A3(net435),
    .S0(net338),
    .S1(net656),
    .X(net652));
 sky130_fd_sc_hd__mux4_1 merge791 (.A0(net435),
    .A1(net858),
    .A2(net962),
    .A3(net445),
    .S0(net212),
    .S1(net798),
    .X(net653));
 sky130_fd_sc_hd__mux4_1 merge792 (.A0(net437),
    .A1(net1109),
    .A2(net962),
    .A3(net556),
    .S0(net445),
    .S1(net976),
    .X(net654));
 sky130_fd_sc_hd__and2_0 merge793 (.A(net226),
    .B(net228),
    .X(net655));
 sky130_fd_sc_hd__dfrbp_2 merge794 (.CLK(clknet_4_10_0_clk),
    .D(net332),
    .RESET_B(net337),
    .Q(net657),
    .Q_N(net656));
 sky130_fd_sc_hd__and2_0 merge795 (.A(net276),
    .B(net259),
    .X(net658));
 sky130_fd_sc_hd__and2_0 merge796 (.A(net591),
    .B(net592),
    .X(net659));
 sky130_fd_sc_hd__and2_1 merge797 (.A(net242),
    .B(net250),
    .X(net660));
 sky130_fd_sc_hd__dfrbp_1 merge798 (.CLK(clknet_4_10_0_clk),
    .D(net652),
    .RESET_B(net654),
    .Q(net662),
    .Q_N(net661));
 sky130_fd_sc_hd__dfrtn_1 merge799 (.CLK_N(clknet_4_0_0_clk),
    .D(net156),
    .RESET_B(net157),
    .Q(net663));
 sky130_fd_sc_hd__dfrtp_4 merge800 (.CLK(clknet_4_2_0_clk),
    .D(net149),
    .RESET_B(net143),
    .Q(net664));
 sky130_fd_sc_hd__dfrtp_1 merge801 (.CLK(clknet_4_10_0_clk),
    .D(net563),
    .RESET_B(net559),
    .Q(net665));
 sky130_fd_sc_hd__dfrtp_1 merge802 (.CLK(clknet_4_9_0_clk),
    .D(net386),
    .RESET_B(net371),
    .Q(net666));
 sky130_fd_sc_hd__and2_0 merge803 (.A(net391),
    .B(net394),
    .X(net667));
 sky130_fd_sc_hd__and2_0 merge804 (.A(net651),
    .B(net633),
    .X(net668));
 sky130_fd_sc_hd__and2_0 merge805 (.A(net300),
    .B(net309),
    .X(net669));
 sky130_fd_sc_hd__and2_0 merge806 (.A(net525),
    .B(net536),
    .X(net670));
 sky130_fd_sc_hd__and2_0 merge807 (.A(net504),
    .B(net505),
    .X(net671));
 sky130_fd_sc_hd__dfsbp_1 merge808 (.CLK(clknet_4_1_0_clk),
    .D(net290),
    .SET_B(net295),
    .Q(net672),
    .Q_N(net950));
 sky130_fd_sc_hd__dfsbp_1 merge809 (.CLK(clknet_4_0_0_clk),
    .D(net173),
    .SET_B(net174),
    .Q(net674),
    .Q_N(net673));
 sky130_fd_sc_hd__and2_0 merge810 (.A(net572),
    .B(net573),
    .X(net675));
 sky130_fd_sc_hd__dfstp_2 merge811 (.CLK(clknet_4_8_0_clk),
    .D(net350),
    .SET_B(net351),
    .Q(net676));
 sky130_fd_sc_hd__dfstp_2 merge812 (.CLK(clknet_4_10_0_clk),
    .D(net458),
    .SET_B(net460),
    .Q(net677));
 sky130_fd_sc_hd__dfstp_1 merge813 (.CLK(clknet_4_14_0_clk),
    .D(net499),
    .SET_B(net480),
    .Q(net678));
 sky130_fd_sc_hd__and2_0 merge814 (.A(net409),
    .B(net412),
    .X(net679));
 sky130_fd_sc_hd__and2_0 merge815 (.A(net430),
    .B(net431),
    .X(net680));
 sky130_fd_sc_hd__dlrbn_2 merge816 (.D(net128),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net124),
    .Q(net682),
    .Q_N(net681));
 sky130_fd_sc_hd__dlrbn_1 merge817 (.D(net611),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net614),
    .Q(net684),
    .Q_N(net683));
 sky130_fd_sc_hd__dlrbp_2 merge818 (.D(net126),
    .GATE(clknet_4_2_0_clk),
    .RESET_B(net123),
    .Q(net686),
    .Q_N(net685));
 sky130_fd_sc_hd__and2_0 merge819 (.A(net585),
    .B(net582),
    .X(net687));
 sky130_fd_sc_hd__dlrbp_1 merge820 (.D(net594),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net607),
    .Q(net689),
    .Q_N(net688));
 sky130_fd_sc_hd__dlrtn_2 merge821 (.D(net278),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net277),
    .Q(net690));
 sky130_fd_sc_hd__dlrtn_1 merge822 (.D(net142),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net145),
    .Q(net917));
 sky130_fd_sc_hd__dlrtn_2 merge823 (.D(net474),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net441),
    .Q(net691));
 sky130_fd_sc_hd__dlrtp_1 merge824 (.D(net161),
    .GATE(clknet_4_0_0_clk),
    .RESET_B(net175),
    .Q(net692));
 sky130_fd_sc_hd__dlrtp_1 merge825 (.D(net229),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net231),
    .Q(net693));
 sky130_fd_sc_hd__dlrtp_1 merge826 (.D(net564),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net675),
    .Q(net694));
 sky130_fd_sc_hd__and2_0 merge827 (.A(net418),
    .B(net317),
    .X(net695));
 sky130_fd_sc_hd__and2_0 merge828 (.A(net539),
    .B(net668),
    .X(net696));
 sky130_fd_sc_hd__and2_4 merge829 (.A(net312),
    .B(net413),
    .X(net697));
 sky130_fd_sc_hd__edfxbp_1 merge830 (.CLK(clknet_4_0_0_clk),
    .D(net180),
    .Q(net183),
    .Q_N(net698));
 sky130_fd_sc_hd__edfxtp_1 merge831 (.CLK(clknet_4_1_0_clk),
    .D(net266),
    .DE(net185),
    .Q(net700));
 sky130_fd_sc_hd__and2_0 merge832 (.A(net510),
    .B(net646),
    .X(net701));
 sky130_fd_sc_hd__and2_0 merge833 (.A(net649),
    .B(net514),
    .X(net702));
 sky130_fd_sc_hd__and2_0 merge834 (.A(net596),
    .B(net629),
    .X(net703));
 sky130_fd_sc_hd__and2_0 merge835 (.A(net397),
    .B(net543),
    .X(net704));
 sky130_fd_sc_hd__and2_0 merge836 (.A(net597),
    .B(net603),
    .X(net705));
 sky130_fd_sc_hd__sdlclkp_1 merge837 (.CLK(clknet_4_9_0_clk),
    .GATE(net352),
    .SCE(net356),
    .GCLK(net706));
 sky130_fd_sc_hd__sdlclkp_2 merge838 (.CLK(clknet_4_13_0_clk),
    .GATE(net621),
    .GCLK(net707));
 sky130_fd_sc_hd__sdlclkp_4 merge839 (.CLK(clknet_4_4_0_clk),
    .GATE(net669),
    .SCE(net297),
    .GCLK(net948));
 sky130_fd_sc_hd__and2_0 merge840 (.A(net520),
    .B(net401),
    .X(net708));
 sky130_fd_sc_hd__dfrbp_1 merge841 (.CLK(clknet_4_4_0_clk),
    .D(net270),
    .RESET_B(net273),
    .Q(net710),
    .Q_N(net709));
 sky130_fd_sc_hd__and2_0 merge842 (.A(net540),
    .B(net634),
    .X(net711));
 sky130_fd_sc_hd__dfrbp_2 merge843 (.CLK(clknet_4_3_0_clk),
    .D(net251),
    .RESET_B(net256),
    .Q(net712),
    .Q_N(net935));
 sky130_fd_sc_hd__and2_0 merge844 (.A(net428),
    .B(net426),
    .X(net713));
 sky130_fd_sc_hd__and2_0 merge845 (.A(net602),
    .B(net628),
    .X(net714));
 sky130_fd_sc_hd__dfrtn_1 merge846 (.CLK_N(clknet_4_15_0_clk),
    .D(net497),
    .RESET_B(net495),
    .Q(net715));
 sky130_fd_sc_hd__and2_0 merge847 (.A(net637),
    .B(net425),
    .X(net716));
 sky130_fd_sc_hd__dfrtp_2 merge848 (.CLK(clknet_4_6_0_clk),
    .D(net704),
    .RESET_B(net374),
    .Q(net717));
 sky130_fd_sc_hd__dfrtp_4 merge849 (.CLK(clknet_4_0_0_clk),
    .D(net158),
    .RESET_B(net159),
    .Q(net718));
 sky130_fd_sc_hd__and2_0 merge850 (.A(net423),
    .B(net420),
    .X(net719));
 sky130_fd_sc_hd__dfrtp_1 merge851 (.CLK(clknet_4_13_0_clk),
    .D(net521),
    .RESET_B(net680),
    .Q(net960));
 sky130_fd_sc_hd__and2_0 merge852 (.A(net383),
    .B(net381),
    .X(net720));
 sky130_fd_sc_hd__and2_0 merge853 (.A(net643),
    .B(net627),
    .X(net721));
 sky130_fd_sc_hd__dfsbp_1 merge854 (.CLK(clknet_4_13_0_clk),
    .D(net516),
    .SET_B(net711),
    .Q(net723),
    .Q_N(net722));
 sky130_fd_sc_hd__dfsbp_1 merge855 (.CLK(clknet_4_12_0_clk),
    .D(net377),
    .SET_B(net491),
    .Q(net725),
    .Q_N(net724));
 sky130_fd_sc_hd__dfstp_1 merge856 (.CLK(clknet_4_4_0_clk),
    .D(net272),
    .SET_B(net658),
    .Q(net726));
 sky130_fd_sc_hd__dfstp_1 merge857 (.CLK(clknet_4_2_0_clk),
    .D(net660),
    .SET_B(net655),
    .Q(net727));
 sky130_fd_sc_hd__dfstp_2 merge858 (.CLK(clknet_4_1_0_clk),
    .D(net257),
    .SET_B(net315),
    .Q(net949));
 sky130_fd_sc_hd__dlrbn_1 merge859 (.D(net616),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net642),
    .Q(net729),
    .Q_N(net728));
 sky130_fd_sc_hd__and2_0 merge860 (.A(net626),
    .B(net617),
    .X(net730));
 sky130_fd_sc_hd__and2_0 merge861 (.A(net623),
    .B(net635),
    .X(net731));
 sky130_fd_sc_hd__dlrbn_1 merge862 (.GATE_N(clknet_4_14_0_clk),
    .RESET_B(net489),
    .Q(net733),
    .Q_N(net490));
 sky130_fd_sc_hd__dlrbp_1 merge863 (.D(net720),
    .GATE(clknet_4_12_0_clk),
    .RESET_B(net379),
    .Q(net735),
    .Q_N(net734));
 sky130_fd_sc_hd__and2_0 merge864 (.A(net620),
    .B(net641),
    .X(net736));
 sky130_fd_sc_hd__dlrbp_1 merge865 (.D(net697),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net376),
    .Q(net738),
    .Q_N(net737));
 sky130_fd_sc_hd__dlrtn_1 merge866 (.D(net622),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net577),
    .Q(net739));
 sky130_fd_sc_hd__dlrtn_2 merge867 (.D(net636),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net387),
    .Q(net740));
 sky130_fd_sc_hd__dlrtn_1 merge868 (.D(net667),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net408),
    .Q(net741));
 sky130_fd_sc_hd__dlrtp_2 merge869 (.GATE(clknet_4_14_0_clk),
    .RESET_B(net705),
    .Q(net742));
 sky130_fd_sc_hd__dlrtp_1 merge870 (.D(net719),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net670),
    .Q(net924));
 sky130_fd_sc_hd__dlrtp_2 merge871 (.D(net671),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net736),
    .Q(net915));
 sky130_fd_sc_hd__edfxbp_1 merge872 (.CLK(clknet_4_12_0_clk),
    .D(net708),
    .DE(net484),
    .Q(net744),
    .Q_N(net743));
 sky130_fd_sc_hd__edfxtp_1 merge873 (.CLK(clknet_4_4_0_clk),
    .D(net405),
    .DE(net713),
    .Q(net745));
 sky130_fd_sc_hd__sdlclkp_1 merge874 (.CLK(clknet_4_15_0_clk),
    .GATE(net731),
    .SCE(net721),
    .GCLK(net916));
 sky130_fd_sc_hd__sdlclkp_2 merge875 (.CLK(clknet_4_13_0_clk),
    .GATE(net701),
    .SCE(net696),
    .GCLK(net746));
 sky130_fd_sc_hd__sdlclkp_4 merge876 (.CLK(clknet_4_15_0_clk),
    .GATE(net702),
    .SCE(net579),
    .GCLK(net747));
 sky130_fd_sc_hd__dfrbp_1 merge877 (.CLK(clknet_4_15_0_clk),
    .D(net659),
    .RESET_B(net714),
    .Q(net749),
    .Q_N(net748));
 sky130_fd_sc_hd__dfrbp_2 merge878 (.CLK(clknet_4_4_0_clk),
    .D(net695),
    .RESET_B(net679),
    .Q(net751),
    .Q_N(net750));
 sky130_fd_sc_hd__dfrtn_1 merge879 (.CLK_N(clknet_4_0_0_clk),
    .D(net165),
    .RESET_B(net298),
    .Q(net752));
 sky130_fd_sc_hd__dfrtp_4 merge880 (.CLK(clknet_4_14_0_clk),
    .D(net503),
    .RESET_B(net586),
    .Q(net753));
 sky130_fd_sc_hd__dfrtp_2 merge881 (.CLK(clknet_4_13_0_clk),
    .D(net502),
    .RESET_B(net716),
    .Q(net954));
 sky130_fd_sc_hd__dfrtp_2 merge882 (.CLK(clknet_4_13_0_clk),
    .D(net417),
    .RESET_B(net589),
    .Q(net754));
 sky130_fd_sc_hd__dfsbp_1 merge883 (.CLK(clknet_4_14_0_clk),
    .D(net605),
    .SET_B(net687),
    .Q(net756),
    .Q_N(net755));
 sky130_fd_sc_hd__dfsbp_2 merge884 (.CLK(clknet_4_5_0_clk),
    .SET_B(net424),
    .Q(net757),
    .Q_N(net429));
 sky130_fd_sc_hd__dfstp_2 merge885 (.CLK(clknet_4_1_0_clk),
    .D(net260),
    .SET_B(net313),
    .Q(net758));
 sky130_fd_sc_hd__dfstp_1 merge886 (.CLK(clknet_4_13_0_clk),
    .D(net730),
    .SET_B(net511),
    .Q(net759));
 sky130_fd_sc_hd__dfstp_1 merge887 (.CLK(clknet_4_14_0_clk),
    .D(net482),
    .SET_B(net703),
    .Q(net760));
 sky130_fd_sc_hd__dlrbn_2 merge888 (.D(net160),
    .GATE_N(clknet_4_0_0_clk),
    .RESET_B(net293),
    .Q(net761),
    .Q_N(net956));
 sky130_fd_sc_hd__dfxbp_2 s889 (.CLK(clknet_4_2_0_clk),
    .D(net127),
    .Q(net763),
    .Q_N(net762));
 sky130_fd_sc_hd__dfxbp_2 s890 (.CLK(clknet_4_4_0_clk),
    .D(net150),
    .Q(net909),
    .Q_N(net764));
 sky130_fd_sc_hd__dfxtp_4 s891 (.CLK(clknet_4_1_0_clk),
    .D(net167),
    .Q(net765));
 sky130_fd_sc_hd__dfxtp_1 s892 (.CLK(clknet_4_0_0_clk),
    .D(net168),
    .Q(net766));
 sky130_fd_sc_hd__dfxtp_1 s893 (.CLK(clknet_4_0_0_clk),
    .D(net184),
    .Q(net940));
 sky130_fd_sc_hd__dlclkp_1 s894 (.CLK(clknet_4_1_0_clk),
    .GATE(net187),
    .GCLK(net925));
 sky130_fd_sc_hd__dlclkp_2 s895 (.CLK(clknet_4_8_0_clk),
    .GATE(net225),
    .GCLK(net767));
 sky130_fd_sc_hd__dlclkp_4 s896 (.CLK(clknet_4_3_0_clk),
    .GATE(net249),
    .GCLK(net768));
 sky130_fd_sc_hd__dlxbn_2 s897 (.D(net263),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net770),
    .Q_N(net769));
 sky130_fd_sc_hd__dlxbn_1 s898 (.D(net265),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net772),
    .Q_N(net771));
 sky130_fd_sc_hd__dlxbp_1 s899 (.D(net267),
    .GATE(clknet_4_6_0_clk),
    .Q(net774),
    .Q_N(net773));
 sky130_fd_sc_hd__dlxtn_4 s900 (.D(net268),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net945));
 sky130_fd_sc_hd__dlxtn_2 s901 (.D(net271),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net775));
 sky130_fd_sc_hd__dlxtn_4 s902 (.D(net274),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net776));
 sky130_fd_sc_hd__dlxtp_1 s903 (.D(net286),
    .GATE(clknet_4_5_0_clk),
    .Q(net777));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s904 (.D(net289),
    .SLEEP_B(clknet_4_6_0_clk),
    .Q(net778));
 sky130_fd_sc_hd__dfxbp_1 s905 (.CLK(clknet_4_4_0_clk),
    .D(net291),
    .Q(net780),
    .Q_N(net779));
 sky130_fd_sc_hd__dfxbp_1 s906 (.CLK(clknet_4_4_0_clk),
    .D(net292),
    .Q(net782),
    .Q_N(net781));
 sky130_fd_sc_hd__dfxtp_1 s907 (.CLK(clknet_4_1_0_clk),
    .D(net301),
    .Q(net783));
 sky130_fd_sc_hd__dfxtp_1 s908 (.CLK(clknet_4_8_0_clk),
    .D(net344),
    .Q(net784));
 sky130_fd_sc_hd__dfxtp_2 s909 (.CLK(clknet_4_8_0_clk),
    .D(net355),
    .Q(net785));
 sky130_fd_sc_hd__dlclkp_1 s910 (.CLK(clknet_4_11_0_clk),
    .GATE(net359),
    .GCLK(net786));
 sky130_fd_sc_hd__dlclkp_2 s911 (.CLK(clknet_4_8_0_clk),
    .GATE(net360),
    .GCLK(net951));
 sky130_fd_sc_hd__dlclkp_4 s912 (.CLK(clknet_4_9_0_clk),
    .GATE(net362),
    .GCLK(net787));
 sky130_fd_sc_hd__dlxbn_1 s913 (.D(net363),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net941),
    .Q_N(net788));
 sky130_fd_sc_hd__dlxbn_1 s914 (.D(net364),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net790),
    .Q_N(net789));
 sky130_fd_sc_hd__dlxbp_1 s915 (.D(net388),
    .GATE(clknet_4_6_0_clk),
    .Q(net792),
    .Q_N(net791));
 sky130_fd_sc_hd__dlxtn_2 s916 (.D(net395),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net793));
 sky130_fd_sc_hd__dlxtn_4 s917 (.D(net398),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net928));
 sky130_fd_sc_hd__dlxtn_1 s918 (.D(net406),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net794));
 sky130_fd_sc_hd__dlxtp_1 s919 (.D(net410),
    .GATE(clknet_4_5_0_clk),
    .Q(net938));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s920 (.D(net411),
    .SLEEP_B(clknet_4_6_0_clk),
    .Q(net795));
 sky130_fd_sc_hd__dfxbp_1 s921 (.CLK(clknet_4_7_0_clk),
    .D(net415),
    .Q(net797),
    .Q_N(net796));
 sky130_fd_sc_hd__dfxbp_1 s922 (.CLK(clknet_4_10_0_clk),
    .D(net452),
    .Q(net799),
    .Q_N(net798));
 sky130_fd_sc_hd__dfxtp_4 s923 (.CLK(clknet_4_11_0_clk),
    .D(net459),
    .Q(net800));
 sky130_fd_sc_hd__dfxtp_1 s924 (.CLK(clknet_4_11_0_clk),
    .D(net465),
    .Q(net801));
 sky130_fd_sc_hd__dfxtp_1 s925 (.CLK(clknet_4_9_0_clk),
    .D(net472),
    .Q(net802));
 sky130_fd_sc_hd__dlclkp_1 s926 (.CLK(clknet_4_11_0_clk),
    .GATE(net475),
    .GCLK(net803));
 sky130_fd_sc_hd__dlclkp_2 s927 (.CLK(clknet_4_14_0_clk),
    .GATE(net481),
    .GCLK(net804));
 sky130_fd_sc_hd__dlclkp_4 s928 (.CLK(clknet_4_12_0_clk),
    .GATE(net483),
    .GCLK(net805));
 sky130_fd_sc_hd__dlxbn_1 s929 (.D(net486),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net807),
    .Q_N(net806));
 sky130_fd_sc_hd__dlxbn_1 s930 (.D(net487),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net907),
    .Q_N(net808));
 sky130_fd_sc_hd__dlxbp_1 s931 (.D(net488),
    .GATE(clknet_4_12_0_clk),
    .Q(net810),
    .Q_N(net809));
 sky130_fd_sc_hd__dlxtn_1 s932 (.D(net494),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net811));
 sky130_fd_sc_hd__dlxtn_1 s933 (.D(net501),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net812));
 sky130_fd_sc_hd__dlxtn_2 s934 (.D(net506),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net813));
 sky130_fd_sc_hd__dlxtp_1 s935 (.D(net509),
    .GATE(clknet_4_7_0_clk),
    .Q(net958));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s936 (.D(net515),
    .SLEEP_B(clknet_4_13_0_clk),
    .Q(net814));
 sky130_fd_sc_hd__dfxbp_1 s937 (.CLK(clknet_4_13_0_clk),
    .D(net519),
    .Q(net816),
    .Q_N(net815));
 sky130_fd_sc_hd__dfxbp_1 s938 (.CLK(clknet_4_7_0_clk),
    .D(net522),
    .Q(net818),
    .Q_N(net817));
 sky130_fd_sc_hd__dfxtp_1 s939 (.CLK(clknet_4_5_0_clk),
    .D(net523),
    .Q(net922));
 sky130_fd_sc_hd__dfxtp_1 s940 (.CLK(clknet_4_7_0_clk),
    .D(net524),
    .Q(net819));
 sky130_fd_sc_hd__dfxtp_1 s941 (.CLK(clknet_4_7_0_clk),
    .D(net527),
    .Q(net820));
 sky130_fd_sc_hd__dlclkp_1 s942 (.CLK(clknet_4_7_0_clk),
    .GATE(net532),
    .GCLK(net821));
 sky130_fd_sc_hd__dlclkp_2 s943 (.CLK(clknet_4_5_0_clk),
    .GATE(net533),
    .GCLK(net822));
 sky130_fd_sc_hd__dlclkp_4 s944 (.CLK(clknet_4_7_0_clk),
    .GATE(net538),
    .GCLK(net823));
 sky130_fd_sc_hd__dlxbn_1 s945 (.D(net562),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net825),
    .Q_N(net824));
 sky130_fd_sc_hd__dlxbn_1 s946 (.D(net565),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net827),
    .Q_N(net826));
 sky130_fd_sc_hd__dlxbp_1 s947 (.D(net566),
    .GATE(clknet_4_11_0_clk),
    .Q(net829),
    .Q_N(net828));
 sky130_fd_sc_hd__dlxtn_2 s948 (.D(net574),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net830));
 sky130_fd_sc_hd__dlxtn_1 s949 (.D(net576),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net831));
 sky130_fd_sc_hd__dlxtn_1 s950 (.D(net578),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net912));
 sky130_fd_sc_hd__dlxtp_1 s951 (.D(net580),
    .GATE(clknet_4_11_0_clk),
    .Q(net832));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s952 (.D(net583),
    .SLEEP_B(clknet_4_11_0_clk),
    .Q(net833));
 sky130_fd_sc_hd__dfxbp_1 s953 (.CLK(clknet_4_14_0_clk),
    .D(net588),
    .Q(net835),
    .Q_N(net834));
 sky130_fd_sc_hd__dfxbp_1 s954 (.CLK(clknet_4_14_0_clk),
    .D(net590),
    .Q(net837),
    .Q_N(net836));
 sky130_fd_sc_hd__dfxtp_1 s955 (.CLK(clknet_4_14_0_clk),
    .D(net593),
    .Q(net838));
 sky130_fd_sc_hd__dfxtp_1 s956 (.CLK(clknet_4_14_0_clk),
    .D(net595),
    .Q(net839));
 sky130_fd_sc_hd__dfxtp_1 s957 (.CLK(clknet_4_14_0_clk),
    .D(net599),
    .Q(net840));
 sky130_fd_sc_hd__dlclkp_1 s958 (.CLK(clknet_4_15_0_clk),
    .GATE(net600),
    .GCLK(net841));
 sky130_fd_sc_hd__dlclkp_2 s959 (.CLK(clknet_4_15_0_clk),
    .GATE(net624),
    .GCLK(net842));
 sky130_fd_sc_hd__dlclkp_4 s960 (.CLK(clknet_4_15_0_clk),
    .GATE(net625),
    .GCLK(net843));
 sky130_fd_sc_hd__dlxbn_1 s961 (.D(net653),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net845),
    .Q_N(net844));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(in0),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(in1),
    .X(net645));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(in10),
    .X(net846));
 sky130_fd_sc_hd__buf_2 input4 (.A(in11),
    .X(net847));
 sky130_fd_sc_hd__buf_8 input5 (.A(in12),
    .X(net848));
 sky130_fd_sc_hd__buf_1 input6 (.A(in13),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(in14),
    .X(net850));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(in15),
    .X(net851));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(in16),
    .X(net852));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(in17),
    .X(net853));
 sky130_fd_sc_hd__buf_2 input11 (.A(in18),
    .X(net854));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(in19),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(in2),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(in20),
    .X(net857));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(in21),
    .X(net858));
 sky130_fd_sc_hd__buf_4 input16 (.A(in22),
    .X(net859));
 sky130_fd_sc_hd__buf_2 input17 (.A(in23),
    .X(net860));
 sky130_fd_sc_hd__buf_2 input18 (.A(in24),
    .X(net861));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(in25),
    .X(net862));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(in26),
    .X(net863));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(in27),
    .X(net864));
 sky130_fd_sc_hd__buf_2 input22 (.A(in28),
    .X(net865));
 sky130_fd_sc_hd__buf_4 input23 (.A(in29),
    .X(net866));
 sky130_fd_sc_hd__buf_2 input24 (.A(in3),
    .X(net867));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(in30),
    .X(net868));
 sky130_fd_sc_hd__buf_4 input26 (.A(in31),
    .X(net869));
 sky130_fd_sc_hd__buf_4 input27 (.A(in32),
    .X(net870));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(in33),
    .X(net871));
 sky130_fd_sc_hd__buf_2 input29 (.A(in34),
    .X(net872));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(in35),
    .X(net873));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(in36),
    .X(net874));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(in37),
    .X(net875));
 sky130_fd_sc_hd__buf_4 input33 (.A(in38),
    .X(net876));
 sky130_fd_sc_hd__buf_2 input34 (.A(in39),
    .X(net877));
 sky130_fd_sc_hd__buf_1 input35 (.A(in4),
    .X(net878));
 sky130_fd_sc_hd__buf_4 input36 (.A(in40),
    .X(net879));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(in41),
    .X(net880));
 sky130_fd_sc_hd__buf_2 input38 (.A(in42),
    .X(net881));
 sky130_fd_sc_hd__buf_2 input39 (.A(in43),
    .X(net882));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(in44),
    .X(net883));
 sky130_fd_sc_hd__buf_2 input41 (.A(in45),
    .X(net884));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(in46),
    .X(net885));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(in47),
    .X(net886));
 sky130_fd_sc_hd__buf_4 input44 (.A(in48),
    .X(net887));
 sky130_fd_sc_hd__clkbuf_4 input45 (.A(in49),
    .X(net888));
 sky130_fd_sc_hd__buf_1 input46 (.A(in5),
    .X(net889));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(in50),
    .X(net890));
 sky130_fd_sc_hd__clkbuf_4 input48 (.A(in51),
    .X(net891));
 sky130_fd_sc_hd__dlymetal6s2s_1 input49 (.A(in52),
    .X(net892));
 sky130_fd_sc_hd__clkbuf_4 input50 (.A(in53),
    .X(net893));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(in54),
    .X(net894));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(in55),
    .X(net895));
 sky130_fd_sc_hd__buf_2 input53 (.A(in56),
    .X(net896));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(in57),
    .X(net897));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(in58),
    .X(net898));
 sky130_fd_sc_hd__clkbuf_4 input56 (.A(in59),
    .X(net899));
 sky130_fd_sc_hd__dlymetal6s2s_1 input57 (.A(in6),
    .X(net900));
 sky130_fd_sc_hd__buf_2 input58 (.A(in60),
    .X(net901));
 sky130_fd_sc_hd__buf_2 input59 (.A(in61),
    .X(net902));
 sky130_fd_sc_hd__buf_4 input60 (.A(in7),
    .X(net903));
 sky130_fd_sc_hd__buf_2 input61 (.A(in8),
    .X(net904));
 sky130_fd_sc_hd__buf_2 input62 (.A(in9),
    .X(net905));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(net906),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net907),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output65 (.A(net908),
    .X(out10));
 sky130_fd_sc_hd__clkbuf_4 output66 (.A(net909),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output67 (.A(net993),
    .X(out14));
 sky130_fd_sc_hd__clkbuf_4 output68 (.A(net911),
    .X(out15));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net912),
    .X(out16));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(clknet_1_0__leaf_net913),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output71 (.A(net914),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output72 (.A(net915),
    .X(out19));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(clknet_1_1__leaf_net916),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output74 (.A(net1009),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output75 (.A(net918),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output76 (.A(net919),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_4 output77 (.A(net920),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output78 (.A(net921),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output79 (.A(net922),
    .X(out25));
 sky130_fd_sc_hd__buf_2 output80 (.A(net923),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output81 (.A(net924),
    .X(out27));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(clknet_1_0__leaf_net925),
    .X(out28));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net926),
    .X(out29));
 sky130_fd_sc_hd__buf_2 output84 (.A(net927),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output85 (.A(net928),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output86 (.A(net1014),
    .X(out31));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(clknet_1_0__leaf_net930),
    .X(out32));
 sky130_fd_sc_hd__buf_2 output88 (.A(net967),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output89 (.A(net1012),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output90 (.A(net933),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_4 output91 (.A(net934),
    .X(out37));
 sky130_fd_sc_hd__buf_2 output92 (.A(net935),
    .X(out38));
 sky130_fd_sc_hd__buf_2 output93 (.A(net971),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_4 output94 (.A(net937),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output95 (.A(net938),
    .X(out41));
 sky130_fd_sc_hd__buf_2 output96 (.A(net1054),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output97 (.A(net940),
    .X(out43));
 sky130_fd_sc_hd__clkbuf_4 output98 (.A(net941),
    .X(out44));
 sky130_fd_sc_hd__buf_2 output99 (.A(net942),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output100 (.A(net943),
    .X(out46));
 sky130_fd_sc_hd__buf_2 output101 (.A(net944),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output102 (.A(net945),
    .X(out48));
 sky130_fd_sc_hd__buf_2 output103 (.A(net946),
    .X(out49));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net963),
    .X(out5));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(clknet_1_0__leaf_net948),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output106 (.A(net949),
    .X(out51));
 sky130_fd_sc_hd__buf_2 output107 (.A(net950),
    .X(out52));
 sky130_fd_sc_hd__clkbuf_1 output108 (.A(clknet_1_1__leaf_net951),
    .X(out53));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(clknet_1_0__leaf_net952),
    .X(out54));
 sky130_fd_sc_hd__clkbuf_1 output110 (.A(clknet_1_0__leaf_net953),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output111 (.A(net954),
    .X(out56));
 sky130_fd_sc_hd__buf_2 output112 (.A(net955),
    .X(out57));
 sky130_fd_sc_hd__buf_2 output113 (.A(net956),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output114 (.A(net965),
    .X(out61));
 sky130_fd_sc_hd__buf_2 output115 (.A(net958),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_4 output116 (.A(net959),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output117 (.A(net960),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_4 fanout118 (.A(net455),
    .X(net961));
 sky130_fd_sc_hd__clkbuf_4 fanout119 (.A(net963),
    .X(net962));
 sky130_fd_sc_hd__clkbuf_4 fanout120 (.A(net947),
    .X(net963));
 sky130_fd_sc_hd__clkbuf_4 fanout121 (.A(net959),
    .X(net964));
 sky130_fd_sc_hd__buf_4 fanout122 (.A(net957),
    .X(net965));
 sky130_fd_sc_hd__clkbuf_4 fanout123 (.A(net340),
    .X(net966));
 sky130_fd_sc_hd__buf_4 fanout124 (.A(net931),
    .X(net967));
 sky130_fd_sc_hd__clkbuf_4 fanout125 (.A(net108),
    .X(net968));
 sky130_fd_sc_hd__buf_2 fanout126 (.A(net970),
    .X(net969));
 sky130_fd_sc_hd__buf_2 fanout127 (.A(net971),
    .X(net970));
 sky130_fd_sc_hd__buf_4 fanout128 (.A(net936),
    .X(net971));
 sky130_fd_sc_hd__clkbuf_4 fanout129 (.A(net210),
    .X(net972));
 sky130_fd_sc_hd__clkbuf_2 fanout130 (.A(net210),
    .X(net973));
 sky130_fd_sc_hd__buf_6 fanout131 (.A(net106),
    .X(net974));
 sky130_fd_sc_hd__clkbuf_4 fanout132 (.A(net208),
    .X(net975));
 sky130_fd_sc_hd__buf_2 fanout133 (.A(net208),
    .X(net976));
 sky130_fd_sc_hd__clkbuf_4 fanout134 (.A(net937),
    .X(net977));
 sky130_fd_sc_hd__clkbuf_4 fanout135 (.A(net979),
    .X(net978));
 sky130_fd_sc_hd__buf_8 fanout136 (.A(net980),
    .X(net979));
 sky130_fd_sc_hd__buf_6 fanout137 (.A(net98),
    .X(net980));
 sky130_fd_sc_hd__buf_8 fanout138 (.A(net32),
    .X(net981));
 sky130_fd_sc_hd__buf_4 fanout139 (.A(net319),
    .X(net982));
 sky130_fd_sc_hd__buf_4 fanout140 (.A(net95),
    .X(net983));
 sky130_fd_sc_hd__clkbuf_2 fanout141 (.A(net95),
    .X(net984));
 sky130_fd_sc_hd__clkbuf_4 fanout142 (.A(net91),
    .X(net985));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout143 (.A(net91),
    .X(net986));
 sky130_fd_sc_hd__buf_8 fanout144 (.A(net24),
    .X(net987));
 sky130_fd_sc_hd__clkbuf_2 fanout145 (.A(net1125),
    .X(net988));
 sky130_fd_sc_hd__buf_8 fanout146 (.A(net84),
    .X(net989));
 sky130_fd_sc_hd__buf_6 fanout147 (.A(net81),
    .X(net990));
 sky130_fd_sc_hd__buf_8 fanout148 (.A(net20),
    .X(net991));
 sky130_fd_sc_hd__buf_8 fanout149 (.A(net993),
    .X(net992));
 sky130_fd_sc_hd__buf_6 fanout150 (.A(net910),
    .X(net993));
 sky130_fd_sc_hd__buf_4 fanout151 (.A(net78),
    .X(net994));
 sky130_fd_sc_hd__clkbuf_2 fanout152 (.A(net78),
    .X(net995));
 sky130_fd_sc_hd__buf_6 fanout153 (.A(net77),
    .X(net996));
 sky130_fd_sc_hd__buf_6 fanout154 (.A(net76),
    .X(net997));
 sky130_fd_sc_hd__clkbuf_4 fanout155 (.A(net88),
    .X(net998));
 sky130_fd_sc_hd__clkbuf_4 fanout156 (.A(net549),
    .X(net999));
 sky130_fd_sc_hd__buf_4 fanout157 (.A(net323),
    .X(net1000));
 sky130_fd_sc_hd__clkbuf_4 fanout158 (.A(net1002),
    .X(net1001));
 sky130_fd_sc_hd__buf_6 fanout159 (.A(net1003),
    .X(net1002));
 sky130_fd_sc_hd__buf_4 fanout160 (.A(net1004),
    .X(net1003));
 sky130_fd_sc_hd__buf_6 fanout161 (.A(net72),
    .X(net1004));
 sky130_fd_sc_hd__clkbuf_4 fanout162 (.A(net778),
    .X(net1005));
 sky130_fd_sc_hd__buf_4 fanout163 (.A(net727),
    .X(net1006));
 sky130_fd_sc_hd__buf_2 fanout164 (.A(net727),
    .X(net1007));
 sky130_fd_sc_hd__buf_4 fanout165 (.A(net693),
    .X(net1008));
 sky130_fd_sc_hd__buf_4 fanout166 (.A(net917),
    .X(net1009));
 sky130_fd_sc_hd__clkbuf_4 fanout167 (.A(net140),
    .X(net1010));
 sky130_fd_sc_hd__clkbuf_4 fanout168 (.A(net1012),
    .X(net1011));
 sky130_fd_sc_hd__clkbuf_4 fanout169 (.A(net932),
    .X(net1012));
 sky130_fd_sc_hd__buf_6 fanout170 (.A(net70),
    .X(net1013));
 sky130_fd_sc_hd__clkbuf_4 fanout171 (.A(net929),
    .X(net1014));
 sky130_fd_sc_hd__buf_2 fanout172 (.A(net929),
    .X(net1015));
 sky130_fd_sc_hd__buf_4 fanout173 (.A(net852),
    .X(net1016));
 sky130_fd_sc_hd__buf_4 fanout174 (.A(net851),
    .X(net1017));
 sky130_fd_sc_hd__clkbuf_8 fanout175 (.A(net850),
    .X(net1018));
 sky130_fd_sc_hd__buf_2 fanout176 (.A(net850),
    .X(net1019));
 sky130_fd_sc_hd__clkbuf_8 fanout177 (.A(net905),
    .X(net1020));
 sky130_fd_sc_hd__clkbuf_4 fanout178 (.A(net904),
    .X(net1021));
 sky130_fd_sc_hd__buf_4 fanout179 (.A(net849),
    .X(net1022));
 sky130_fd_sc_hd__clkbuf_4 fanout180 (.A(net900),
    .X(net1023));
 sky130_fd_sc_hd__buf_2 fanout181 (.A(net1026),
    .X(net1024));
 sky130_fd_sc_hd__buf_2 fanout182 (.A(net1026),
    .X(net1025));
 sky130_fd_sc_hd__buf_4 fanout183 (.A(net895),
    .X(net1026));
 sky130_fd_sc_hd__buf_8 fanout184 (.A(net1028),
    .X(net1027));
 sky130_fd_sc_hd__buf_12 fanout185 (.A(net848),
    .X(net1028));
 sky130_fd_sc_hd__buf_4 fanout186 (.A(net892),
    .X(net1029));
 sky130_fd_sc_hd__buf_2 fanout187 (.A(net892),
    .X(net1030));
 sky130_fd_sc_hd__buf_4 fanout188 (.A(net889),
    .X(net1031));
 sky130_fd_sc_hd__buf_4 fanout189 (.A(net885),
    .X(net1032));
 sky130_fd_sc_hd__clkbuf_4 fanout190 (.A(net847),
    .X(net1033));
 sky130_fd_sc_hd__clkbuf_4 fanout191 (.A(net878),
    .X(net1034));
 sky130_fd_sc_hd__buf_4 fanout192 (.A(net875),
    .X(net1035));
 sky130_fd_sc_hd__clkbuf_4 fanout193 (.A(net846),
    .X(net1036));
 sky130_fd_sc_hd__buf_4 fanout194 (.A(net868),
    .X(net1037));
 sky130_fd_sc_hd__buf_12 fanout195 (.A(net867),
    .X(net1038));
 sky130_fd_sc_hd__clkbuf_8 fanout196 (.A(net645),
    .X(net1039));
 sky130_fd_sc_hd__buf_12 fanout197 (.A(net857),
    .X(net1040));
 sky130_fd_sc_hd__buf_8 fanout198 (.A(net856),
    .X(net1041));
 sky130_fd_sc_hd__buf_4 fanout199 (.A(net855),
    .X(net1042));
 sky130_fd_sc_hd__clkbuf_4 fanout200 (.A(net1044),
    .X(net1043));
 sky130_fd_sc_hd__buf_4 fanout201 (.A(net854),
    .X(net1044));
 sky130_fd_sc_hd__clkbuf_4 fanout202 (.A(net853),
    .X(net1045));
 sky130_fd_sc_hd__buf_2 fanout203 (.A(net608),
    .X(net1046));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net843 (.A(net843),
    .X(clknet_0_net843));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net843 (.A(clknet_0_net843),
    .X(clknet_1_0__leaf_net843));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net843 (.A(clknet_0_net843),
    .X(clknet_1_1__leaf_net843));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net916 (.A(net916),
    .X(clknet_0_net916));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net916 (.A(clknet_0_net916),
    .X(clknet_1_0__leaf_net916));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net916 (.A(clknet_0_net916),
    .X(clknet_1_1__leaf_net916));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net746 (.A(net746),
    .X(clknet_0_net746));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net746 (.A(clknet_0_net746),
    .X(clknet_1_0__leaf_net746));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net746 (.A(clknet_0_net746),
    .X(clknet_1_1__leaf_net746));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net747 (.A(net747),
    .X(clknet_0_net747));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net747 (.A(clknet_0_net747),
    .X(clknet_1_0__leaf_net747));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net747 (.A(clknet_0_net747),
    .X(clknet_1_1__leaf_net747));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net821 (.A(net821),
    .X(clknet_0_net821));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net821 (.A(clknet_0_net821),
    .X(clknet_1_0__leaf_net821));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net821 (.A(clknet_0_net821),
    .X(clknet_1_1__leaf_net821));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net542 (.A(net542),
    .X(clknet_0_net542));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net542 (.A(clknet_0_net542),
    .X(clknet_1_0__leaf_net542));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net542 (.A(clknet_0_net542),
    .X(clknet_1_1__leaf_net542));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net842 (.A(net842),
    .X(clknet_0_net842));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net842 (.A(clknet_0_net842),
    .X(clknet_1_0__leaf_net842));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net842 (.A(clknet_0_net842),
    .X(clknet_1_1__leaf_net842));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net841 (.A(net841),
    .X(clknet_0_net841));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net841 (.A(clknet_0_net841),
    .X(clknet_1_0__leaf_net841));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net841 (.A(clknet_0_net841),
    .X(clknet_1_1__leaf_net841));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net604 (.A(net604),
    .X(clknet_0_net604));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net604 (.A(clknet_0_net604),
    .X(clknet_1_0__leaf_net604));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net604 (.A(clknet_0_net604),
    .X(clknet_1_1__leaf_net604));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net742 (.A(net742),
    .X(clknet_0_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net742 (.A(clknet_0_net742),
    .X(clknet_1_0__leaf_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net742 (.A(clknet_0_net742),
    .X(clknet_1_1__leaf_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net823 (.A(net823),
    .X(clknet_0_net823));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net823 (.A(clknet_0_net823),
    .X(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net823 (.A(clknet_0_net823),
    .X(clknet_1_1__leaf_net823));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net822 (.A(net822),
    .X(clknet_0_net822));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net822 (.A(clknet_0_net822),
    .X(clknet_1_0__leaf_net822));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net822 (.A(clknet_0_net822),
    .X(clknet_1_1__leaf_net822));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net537 (.A(net537),
    .X(clknet_0_net537));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net537 (.A(clknet_0_net537),
    .X(clknet_1_0__leaf_net537));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net537 (.A(clknet_0_net537),
    .X(clknet_1_1__leaf_net537));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net805 (.A(net805),
    .X(clknet_0_net805));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net805 (.A(clknet_0_net805),
    .X(clknet_1_0__leaf_net805));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net805 (.A(clknet_0_net805),
    .X(clknet_1_1__leaf_net805));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net534 (.A(net534),
    .X(clknet_0_net534));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net534 (.A(clknet_0_net534),
    .X(clknet_1_0__leaf_net534));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net534 (.A(clknet_0_net534),
    .X(clknet_1_1__leaf_net534));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net485 (.A(net485),
    .X(clknet_0_net485));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net485 (.A(clknet_0_net485),
    .X(clknet_1_0__leaf_net485));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net485 (.A(clknet_0_net485),
    .X(clknet_1_1__leaf_net485));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net804 (.A(net804),
    .X(clknet_0_net804));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net804 (.A(clknet_0_net804),
    .X(clknet_1_0__leaf_net804));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net804 (.A(clknet_0_net804),
    .X(clknet_1_1__leaf_net804));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net618 (.A(net618),
    .X(clknet_0_net618));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net618 (.A(clknet_0_net618),
    .X(clknet_1_0__leaf_net618));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net618 (.A(clknet_0_net618),
    .X(clknet_1_1__leaf_net618));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net803 (.A(net803),
    .X(clknet_0_net803));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net803 (.A(clknet_0_net803),
    .X(clknet_1_0__leaf_net803));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net803 (.A(clknet_0_net803),
    .X(clknet_1_1__leaf_net803));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net498 (.A(net498),
    .X(clknet_0_net498));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net498 (.A(clknet_0_net498),
    .X(clknet_1_0__leaf_net498));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net498 (.A(clknet_0_net498),
    .X(clknet_1_1__leaf_net498));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net477 (.A(net477),
    .X(clknet_0_net477));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net477 (.A(clknet_0_net477),
    .X(clknet_1_0__leaf_net477));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net477 (.A(clknet_0_net477),
    .X(clknet_1_1__leaf_net477));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net581 (.A(net581),
    .X(clknet_0_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net581 (.A(clknet_0_net581),
    .X(clknet_1_0__leaf_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net581 (.A(clknet_0_net581),
    .X(clknet_1_1__leaf_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net575 (.A(net575),
    .X(clknet_0_net575));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net575 (.A(clknet_0_net575),
    .X(clknet_1_0__leaf_net575));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net575 (.A(clknet_0_net575),
    .X(clknet_1_1__leaf_net575));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net568 (.A(net568),
    .X(clknet_0_net568));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net568 (.A(clknet_0_net568),
    .X(clknet_1_0__leaf_net568));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net568 (.A(clknet_0_net568),
    .X(clknet_1_1__leaf_net568));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net787 (.A(net787),
    .X(clknet_0_net787));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net787 (.A(clknet_0_net787),
    .X(clknet_1_0__leaf_net787));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net787 (.A(clknet_0_net787),
    .X(clknet_1_1__leaf_net787));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net380 (.A(net380),
    .X(clknet_0_net380));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net380 (.A(clknet_0_net380),
    .X(clknet_1_0__leaf_net380));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net380 (.A(clknet_0_net380),
    .X(clknet_1_1__leaf_net380));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net496 (.A(net496),
    .X(clknet_0_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net496 (.A(clknet_0_net496),
    .X(clknet_1_0__leaf_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net496 (.A(clknet_0_net496),
    .X(clknet_1_1__leaf_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net479 (.A(net479),
    .X(clknet_0_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net479 (.A(clknet_0_net479),
    .X(clknet_1_0__leaf_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net479 (.A(clknet_0_net479),
    .X(clknet_1_1__leaf_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net400 (.A(net400),
    .X(clknet_0_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net400 (.A(clknet_0_net400),
    .X(clknet_1_0__leaf_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net400 (.A(clknet_0_net400),
    .X(clknet_1_1__leaf_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net507 (.A(net507),
    .X(clknet_0_net507));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net507 (.A(clknet_0_net507),
    .X(clknet_1_0__leaf_net507));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net507 (.A(clknet_0_net507),
    .X(clknet_1_1__leaf_net507));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net399 (.A(net399),
    .X(clknet_0_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_0__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_1__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net372 (.A(net372),
    .X(clknet_0_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_0__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_1__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net951 (.A(net951),
    .X(clknet_0_net951));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net951 (.A(clknet_0_net951),
    .X(clknet_1_0__leaf_net951));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net951 (.A(clknet_0_net951),
    .X(clknet_1_1__leaf_net951));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net361 (.A(net361),
    .X(clknet_0_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net361 (.A(clknet_0_net361),
    .X(clknet_1_0__leaf_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net361 (.A(clknet_0_net361),
    .X(clknet_1_1__leaf_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net786 (.A(net786),
    .X(clknet_0_net786));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net786 (.A(clknet_0_net786),
    .X(clknet_1_0__leaf_net786));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net786 (.A(clknet_0_net786),
    .X(clknet_1_1__leaf_net786));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net569 (.A(net569),
    .X(clknet_0_net569));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net569 (.A(clknet_0_net569),
    .X(clknet_1_0__leaf_net569));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net569 (.A(clknet_0_net569),
    .X(clknet_1_1__leaf_net569));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net567 (.A(net567),
    .X(clknet_0_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net567 (.A(clknet_0_net567),
    .X(clknet_1_0__leaf_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net567 (.A(clknet_0_net567),
    .X(clknet_1_1__leaf_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net768 (.A(net768),
    .X(clknet_0_net768));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net768 (.A(clknet_0_net768),
    .X(clknet_1_0__leaf_net768));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net768 (.A(clknet_0_net768),
    .X(clknet_1_1__leaf_net768));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net389 (.A(net389),
    .X(clknet_0_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_0__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_1__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net269 (.A(net269),
    .X(clknet_0_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net269 (.A(clknet_0_net269),
    .X(clknet_1_0__leaf_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net269 (.A(clknet_0_net269),
    .X(clknet_1_1__leaf_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net264 (.A(net264),
    .X(clknet_0_net264));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net264 (.A(clknet_0_net264),
    .X(clknet_1_0__leaf_net264));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net264 (.A(clknet_0_net264),
    .X(clknet_1_1__leaf_net264));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net254 (.A(net254),
    .X(clknet_0_net254));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net254 (.A(clknet_0_net254),
    .X(clknet_1_0__leaf_net254));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net254 (.A(clknet_0_net254),
    .X(clknet_1_1__leaf_net254));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net767 (.A(net767),
    .X(clknet_0_net767));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net767 (.A(clknet_0_net767),
    .X(clknet_1_0__leaf_net767));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net767 (.A(clknet_0_net767),
    .X(clknet_1_1__leaf_net767));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net396 (.A(net396),
    .X(clknet_0_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_0__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_1__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net913 (.A(net913),
    .X(clknet_0_net913));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net913 (.A(clknet_0_net913),
    .X(clknet_1_0__leaf_net913));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net913 (.A(clknet_0_net913),
    .X(clknet_1_1__leaf_net913));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net378 (.A(net378),
    .X(clknet_0_net378));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net378 (.A(clknet_0_net378),
    .X(clknet_1_0__leaf_net378));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net378 (.A(clknet_0_net378),
    .X(clknet_1_1__leaf_net378));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net365 (.A(net365),
    .X(clknet_0_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net365 (.A(clknet_0_net365),
    .X(clknet_1_0__leaf_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net365 (.A(clknet_0_net365),
    .X(clknet_1_1__leaf_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net275 (.A(net275),
    .X(clknet_0_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net275 (.A(clknet_0_net275),
    .X(clknet_1_0__leaf_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net275 (.A(clknet_0_net275),
    .X(clknet_1_1__leaf_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net230 (.A(net230),
    .X(clknet_0_net230));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net230 (.A(clknet_0_net230),
    .X(clknet_1_0__leaf_net230));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net230 (.A(clknet_0_net230),
    .X(clknet_1_1__leaf_net230));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net706 (.A(net706),
    .X(clknet_0_net706));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net706 (.A(clknet_0_net706),
    .X(clknet_1_0__leaf_net706));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net706 (.A(clknet_0_net706),
    .X(clknet_1_1__leaf_net706));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net570 (.A(net570),
    .X(clknet_0_net570));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net570 (.A(clknet_0_net570),
    .X(clknet_1_0__leaf_net570));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net570 (.A(clknet_0_net570),
    .X(clknet_1_1__leaf_net570));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net392 (.A(net392),
    .X(clknet_0_net392));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net392 (.A(clknet_0_net392),
    .X(clknet_1_0__leaf_net392));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net392 (.A(clknet_0_net392),
    .X(clknet_1_1__leaf_net392));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net343 (.A(net343),
    .X(clknet_0_net343));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net343 (.A(clknet_0_net343),
    .X(clknet_1_0__leaf_net343));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net343 (.A(clknet_0_net343),
    .X(clknet_1_1__leaf_net343));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net366 (.A(net366),
    .X(clknet_0_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net366 (.A(clknet_0_net366),
    .X(clknet_1_0__leaf_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net366 (.A(clknet_0_net366),
    .X(clknet_1_1__leaf_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net354 (.A(net354),
    .X(clknet_0_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net354 (.A(clknet_0_net354),
    .X(clknet_1_0__leaf_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net354 (.A(clknet_0_net354),
    .X(clknet_1_1__leaf_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net349 (.A(net349),
    .X(clknet_0_net349));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net349 (.A(clknet_0_net349),
    .X(clknet_1_0__leaf_net349));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net349 (.A(clknet_0_net349),
    .X(clknet_1_1__leaf_net349));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net233 (.A(net233),
    .X(clknet_0_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net233 (.A(clknet_0_net233),
    .X(clknet_1_0__leaf_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net233 (.A(clknet_0_net233),
    .X(clknet_1_1__leaf_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net232 (.A(net232),
    .X(clknet_0_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net232 (.A(clknet_0_net232),
    .X(clknet_1_0__leaf_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net232 (.A(clknet_0_net232),
    .X(clknet_1_1__leaf_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net952 (.A(net952),
    .X(clknet_0_net952));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net952 (.A(clknet_0_net952),
    .X(clknet_1_0__leaf_net952));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net952 (.A(clknet_0_net952),
    .X(clknet_1_1__leaf_net952));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net280 (.A(net280),
    .X(clknet_0_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net280 (.A(clknet_0_net280),
    .X(clknet_1_0__leaf_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net280 (.A(clknet_0_net280),
    .X(clknet_1_1__leaf_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net925 (.A(net925),
    .X(clknet_0_net925));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net925 (.A(clknet_0_net925),
    .X(clknet_1_0__leaf_net925));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net925 (.A(clknet_0_net925),
    .X(clknet_1_1__leaf_net925));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net953 (.A(net953),
    .X(clknet_0_net953));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net953 (.A(clknet_0_net953),
    .X(clknet_1_0__leaf_net953));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net953 (.A(clknet_0_net953),
    .X(clknet_1_1__leaf_net953));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net316 (.A(net316),
    .X(clknet_0_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net316 (.A(clknet_0_net316),
    .X(clknet_1_0__leaf_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net316 (.A(clknet_0_net316),
    .X(clknet_1_1__leaf_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net948 (.A(net948),
    .X(clknet_0_net948));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net948 (.A(clknet_0_net948),
    .X(clknet_1_0__leaf_net948));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net948 (.A(clknet_0_net948),
    .X(clknet_1_1__leaf_net948));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net299 (.A(net299),
    .X(clknet_0_net299));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net299 (.A(clknet_0_net299),
    .X(clknet_1_0__leaf_net299));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net299 (.A(clknet_0_net299),
    .X(clknet_1_1__leaf_net299));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net308 (.A(net308),
    .X(clknet_0_net308));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net308 (.A(clknet_0_net308),
    .X(clknet_1_0__leaf_net308));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net308 (.A(clknet_0_net308),
    .X(clknet_1_1__leaf_net308));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net188 (.A(net188),
    .X(clknet_0_net188));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net188 (.A(clknet_0_net188),
    .X(clknet_1_0__leaf_net188));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net188 (.A(clknet_0_net188),
    .X(clknet_1_1__leaf_net188));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net189 (.A(net189),
    .X(clknet_0_net189));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net189 (.A(clknet_0_net189),
    .X(clknet_1_0__leaf_net189));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net189 (.A(clknet_0_net189),
    .X(clknet_1_1__leaf_net189));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net177 (.A(net177),
    .X(clknet_0_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net177 (.A(clknet_0_net177),
    .X(clknet_1_0__leaf_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net177 (.A(clknet_0_net177),
    .X(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net178 (.A(net178),
    .X(clknet_0_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net178 (.A(clknet_0_net178),
    .X(clknet_1_0__leaf_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net178 (.A(clknet_0_net178),
    .X(clknet_1_1__leaf_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net930 (.A(net930),
    .X(clknet_0_net930));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net930 (.A(clknet_0_net930),
    .X(clknet_1_0__leaf_net930));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net930 (.A(clknet_0_net930),
    .X(clknet_1_1__leaf_net930));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net182 (.A(net182),
    .X(clknet_0_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net182 (.A(clknet_0_net182),
    .X(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net182 (.A(clknet_0_net182),
    .X(clknet_1_1__leaf_net182));
 sky130_fd_sc_hd__mux4_1 clone1 (.A0(net101),
    .A1(net85),
    .A2(net877),
    .A3(net865),
    .S0(net978),
    .S1(net80),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net81),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net81),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net98),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net939),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net1051),
    .X(net1052));
 sky130_fd_sc_hd__clkbuf_1 rebuffer7 (.A(net1052),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net1053),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net42),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net1055),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net94),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net84),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net1073),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net1059),
    .X(net1060));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer15 (.A(net3),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net105),
    .X(net1062));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer17 (.A(net1062),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net1063),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net105),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net1065),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net1066),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net20),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net285),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net1128),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net1070),
    .X(net1071));
 sky130_fd_sc_hd__clkbuf_1 rebuffer26 (.A(net1070),
    .X(net1072));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer27 (.A(net3),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(net1076),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net1074),
    .X(net1075));
 sky130_fd_sc_hd__and3_1 clone30 (.A(net2),
    .B(net1107),
    .C(net1025),
    .X(net1076));
 sky130_fd_sc_hd__clkbuf_1 clone31 (.A(net1078),
    .X(net1077));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer32 (.A(net24),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(net44),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(net1079),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer35 (.A(net55),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer36 (.A(net1083),
    .X(net1082));
 sky130_fd_sc_hd__or4bb_1 clone37 (.A(net1105),
    .B(net85),
    .C_N(net994),
    .D_N(net983),
    .X(net1083));
 sky130_fd_sc_hd__clkbuf_1 clone38 (.A(net20),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer39 (.A(net37),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer40 (.A(net22),
    .X(net1086));
 sky130_fd_sc_hd__clkbuf_1 clone41 (.A(net32),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer42 (.A(net32),
    .X(net1088));
 sky130_fd_sc_hd__clkbuf_1 clone43 (.A(net848),
    .X(net1089));
 sky130_fd_sc_hd__clkbuf_1 clone44 (.A(net856),
    .X(net1090));
 sky130_fd_sc_hd__clkbuf_1 clone45 (.A(net1028),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net784),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net765),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net798),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net828),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net810),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net557),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net335),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net545),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net735),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net820),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net928),
    .X(net1102));
 sky130_fd_sc_hd__clkbuf_1 fanout1 (.A(net978),
    .X(net1103));
 sky130_fd_sc_hd__buf_6 fanout2 (.A(net983),
    .X(net1104));
 sky130_fd_sc_hd__clkbuf_1 fanout3 (.A(net985),
    .X(net1105));
 sky130_fd_sc_hd__buf_4 fanout4 (.A(net994),
    .X(net1106));
 sky130_fd_sc_hd__clkbuf_1 fanout5 (.A(net5),
    .X(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S0 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_X (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A1 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_X (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A3 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A1 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_B1 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A0 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A1 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_SCD (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_C (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A1 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_X (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_X (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A3 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A0 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_C1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A0 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_X (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_S0 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A0 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_C_N (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_C (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_X (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S0 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A0 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_D1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_X (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_S0 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A0 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A3 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_S1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_X (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A0 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_RESET_B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_D1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_D1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_X (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A3 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_D1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_C1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A0 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_X (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_X (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A0 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_X (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_SCE (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_X (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A3 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_C1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_X (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_X (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_S0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A3 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_X (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A0 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A0 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_X (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A0 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_RESET_B (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_X (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A3 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A3 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_S1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_S0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_S1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_C1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_C1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A3 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_Q_N (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_S0 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_X (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A0 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S0 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A3 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_SET_B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A0 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_Q (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_B (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_D_N (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_X (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_B (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A0 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A0 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_X (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_D1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_C1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_X (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A0 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_S0 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A3 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_S0 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_RESET_B (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_X (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_Q (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_X (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A3 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_C (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_C (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_X (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A0 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_X (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A0 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_B (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_X (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A3 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A3 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_S0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A3 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_X (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A3 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_SCE (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_X (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A0 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_C (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_C (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_X (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A3 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_X (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_D (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_C (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_X (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_SCD (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_RESET_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_X (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A0 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A3 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_SCE (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_X (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_X (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A3 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_X (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A0 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A3 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_C (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_X (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_SCD (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A0 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_S0 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_X (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A0 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_D1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A2 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A3 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_X (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A3 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_S0 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_C1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_X (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A0 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_B (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_X (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A3 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A3 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_Q_N (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A2 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A3 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_X (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A2 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S0 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A1 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_X (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_S0 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_C1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S0 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_S0 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_D1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_Q_N (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S0 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A0 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_Q (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_C1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_X (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_B1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_Q_N (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer32_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_X (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A3 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_Q (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A0 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A0 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S0 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A3 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A3 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A3 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_X (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_B1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_X (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_X (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_C1 (.DIODE(net1130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_X (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A2 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A0 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_D (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_C (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_C (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_D_N (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A1 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_A3 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A0 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_X (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S0 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A0 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A0 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_X (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_S0 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_X (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A0 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A3 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_D1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S0 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A0 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A0 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_X (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A0 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A3 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A2 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_X (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A0 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_X (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A3 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_S0 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_X (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_X (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A3 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A3 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A3 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A3 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A3 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_X (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A3 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A0 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A2 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_B (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_X (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A2 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A2 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_C (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_C (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_X (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A3 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A0 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_S0 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_X (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_S1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_X (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_S0 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_S1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_D1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_RESET_B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_D (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_C1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_X (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S0 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A2 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A2 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_X (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_X (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A3 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A3 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_S0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_RESET_B (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A2 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_C1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_SCD (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_Q_N (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold52_A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A3 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A2 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_Q (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A2 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A2 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A2 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_S0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_X (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_S0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A3 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_C_N (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_Q_N (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A2 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_D (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_B1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_Q (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_X (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A0 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A0 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_X (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net343_A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_X (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_Q (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A0 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_S1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A0 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_SET_B (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_B1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_X (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A0 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_S1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_D1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_X (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net349_A (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_X (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A3 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_Q_N (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A0 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A0 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_Q (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_D1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_X (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_S0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_S1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A0 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_D (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A2 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_X (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A0 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_Q (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A3 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_X (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_A3 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_X (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A3 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_C1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_X (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_D (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_X (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_X (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A1 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_SCD (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_D (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_X (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A0 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A3 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A2 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_X (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A0 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A0 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A3 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_RESET_B (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_X (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A0 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_B (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_C (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_X (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A0 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A2 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_S0 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A3 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A3 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_S1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_X (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A3 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A0 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A1 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A2 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A1 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S1 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A0 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_X (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A0 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A0 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A0 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_D (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_X (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A0 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_B1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_X (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S0 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A0 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_B1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_RESET_B (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_D_N (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_X (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A0 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A3 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A1 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_SCE (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_X (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A3 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_C (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_SCE (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_Q_N (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A0 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A0 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_Q (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A2 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A2 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_X (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A1 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A2 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A0 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S0 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A1 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_RESET_B (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_X (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A0 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A1 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A1 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A1 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_X (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A0 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A0 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A3 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_X (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A2 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A3 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A0 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A2 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A3 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_B1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_X (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A3 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S0 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_D1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_X (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S0 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_Q_N (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A0 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_B (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_Q (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A0 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A0 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A3 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_Q (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A3 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A1 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_Q_N (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A0 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_X (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout5_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_X (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A0 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_S0 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A3 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_S1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_C (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_C (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_X (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A0 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_X (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A0 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_S1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A2 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_X (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A0 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_S0 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A2 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A2 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A2 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_X (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A0 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A2 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A2 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_X (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net568_A (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_X (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net569_A (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_X (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A1 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A1 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_X (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_SCE (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_X (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_RESET_B (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_X (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_D_N (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_X (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_D_N (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A2 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_X (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_X (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_Q (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_S1 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_D_N (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S0 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_C1 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A2 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S1 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_Q (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_S1 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S0 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A2 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_D1 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_S1 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_D1 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A3 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_C1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_X (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_RESET_B (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_X (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_Q (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A3 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A3 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S0 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_D1 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_D1 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_Q_N (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_S1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_S1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_S1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_D1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_S1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_Q (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S0 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_D1 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S0 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_B1 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_D1 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S0 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_C1 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A0 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_D (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_D1 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A3 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A2 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S0 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_Q (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_S0 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_S1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S0 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_Q (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_D1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_D1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A3 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_S1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_D_N (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_S1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_C (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_X (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_S0 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_C1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A0 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_X (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_Q (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S0 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A3 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A3 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_S1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_S0 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_B (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A3 (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_B (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A0 (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_X (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_Q (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S0 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A2 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_Q (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A3 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S1 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S1 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A3 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S1 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge848_Q (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A3 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_S0 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A2 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_Q (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S1 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_S1 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S1 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S0 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_C1 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_S1 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_Q_N (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S0 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_B1 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A1 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A0 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A3 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_X (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_Q_N (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S1 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_D1 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_Q (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S0 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_Q (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_S0 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A2 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_S0 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_S0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_X (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_Q (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A2 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S1 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S0 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_Q (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A3 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A3 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S0 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A3 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge877_Q_N (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S1 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S0 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_C1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_S0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_D1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_B (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_X (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_Q (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S0 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_S0 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_S0 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_S0 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_Q (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S0 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S0 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge885_Q (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A3 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_S1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_S1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_S1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge886_Q (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S0 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S0 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A3 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge887_Q (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A2 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A3 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S0 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S0 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_Q_N (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S0 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_S1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_Q (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S0 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S0 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_D1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_Q_N (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S0 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S0 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S1 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold47_A (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_Q (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_S0 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_S1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_S1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_S1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_S1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_S1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_S0 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_S1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A1 (.DIODE(net1129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_B (.DIODE(net1129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_C (.DIODE(net1129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A0 (.DIODE(net1129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net1129));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_Q (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A3 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S0 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S0 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_Q_N (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A3 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_Q (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A3 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S0 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_Q (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S0 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S0 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_S0 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_Q (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_S1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S0 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_S1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_Q (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_S0 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S0 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_S1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_Q (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S1 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S1 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S0 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_Q (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A3 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_S0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_Q_N (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S0 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S0 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_X (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_Q (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S0 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S0 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S0 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_Q (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A3 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A3 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_Q (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S0 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_S1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_D1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_X (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_S0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone1_S1 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A0 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A2 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A1 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A1 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_S1 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A2 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_Q (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S0 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_SCE (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_SCE (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_Q (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A3 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_S0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_Q_N (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S0 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_S0 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_S1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer3_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_A (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A3 (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_X (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold50_A (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_Q (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_Q (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S0 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_S1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_D1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_C (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_D1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A3 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_X (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_s945_Q (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_s946_Q (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_s948_Q (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A3 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A2 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S0 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S0 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_S1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_S0 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_s951_Q (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_S1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_S1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_s952_Q (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer12_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone37_B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone1_A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_S0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_SCD (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A1 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A2 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A0 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B1 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A1 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_C (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A0 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_C (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_X (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_X (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_X (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A1 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_C1 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_B (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A2 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_X (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_S0 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A0 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_D1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A2 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_D (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone43_A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S0 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A3 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A0 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A2 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A1 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone44_A (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A3 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A0 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A3 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_S0 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A2 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_B1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_C1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_SCD (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A0 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S0 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A1 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A3 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_D1 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S0 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A0 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A2 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_A1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A0 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A2 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_A1 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A1 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_B (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A1 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A0 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A0 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A1 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A2 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_B1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A0 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_S0 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A2 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A1 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone1_A3 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A3 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A3 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_S0 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_SCE (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_C1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_D1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_D_N (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_C (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A0 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A0 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A2 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A2 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_B1 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_C1 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S0 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A1 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_D_N (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_B (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A2 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A2 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A0 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A2 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_C (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_S0 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A1 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A0 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_D_N (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_B1 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_X (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A3 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A0 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_C_N (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_C (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_A1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_B (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_A1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A0 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A0 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A1 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A2 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A0 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A3 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_RESET_B (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_S0 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_C1 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A1 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A1 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone1_A2 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_A2 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A2 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_C (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_C (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A1 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S0 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A2 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A3 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A1 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A0 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_D (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A2 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A3 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_C (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A2 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_S0 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_X (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_B (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_A0 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_C_N (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A0 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A2 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_C_N (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_A1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S0 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A0 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_D1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A0 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A0 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A3 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_S0 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S0 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_C1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_C1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_X (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A3 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A0 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A2 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_A (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_C (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A3 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_B1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A0 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A2 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A2 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A0 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A2 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A3 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_X (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_C1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S0 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A3 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_X (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A3 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A0 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_RESET_B (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A2 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A0 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A0 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_D1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_X (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A0 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A0 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A2 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_C (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_A (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_D1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A3 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_D1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_X (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A0 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A3 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_C_N (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A0 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_C (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A3 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_S0 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A0 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_X (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_D1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_C_N (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A2 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_D1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_X (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_Q (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S0 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_S0 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S0 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A2 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_S0 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_C (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_X (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_Q (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A3 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S1 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_Q (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_Q (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A2 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A0 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A3 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A3 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S0 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_X (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A0 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A3 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_RESET_B (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_Q (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S0 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A2 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_C1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_Q (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A3 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A3 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S0 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A2 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A2 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A2 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A3 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A2 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_X (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_A2 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A3 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_D1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_B1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_S0 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_C1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_X (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold56_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_Q (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_S0 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S0 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A0 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S0 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_X (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A2 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_Q (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_X (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_Q_N (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_S1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_S0 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A3 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_X (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_Q (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_S1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A2 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_A3 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A2 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_S1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_C (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_X (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A3 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_X (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_Q (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_S1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_S1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_S1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A0 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_X (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_Q (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_S1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_S0 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_S1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_S1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_Q_N (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S1 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge888_Q_N (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S0 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_C1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A2 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_X (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_s935_Q (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_S1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S0 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S0 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S0 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_S0 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_X (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_X (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_S0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_SET_B (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_RESET_B (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_B1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_S0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_C1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_D (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_SCD (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_X (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_SCE (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_SCD (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_SCD (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_X (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_X (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A0 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A3 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A3 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A0 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A3 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A3 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A3 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_SET_B (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A2 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_X (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A3 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A0 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A3 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_S1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_SCD (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A2 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_S1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A2 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A3 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_X (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A0 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A3 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A3 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_X (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S0 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_S0 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A2 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_X (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_C_N (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A3 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_S0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A3 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_B1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_X (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A2 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_SET_B (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_B1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_C1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_B1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_X (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A3 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A3 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A3 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_X (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_C1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A3 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A3 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_C_N (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_C1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A2 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_C (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A3 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A3 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_X (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A0 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A0 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_X (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_B1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_S0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_D1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_D_N (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A2 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A3 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A2 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A3 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_C (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A0 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A2 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_C1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_C (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_B1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_X (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_S1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_D1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_RESET_B (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_SCE (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_X (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A0 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A0 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A3 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_B1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_B1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A3 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A0 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A3 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_B1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_X (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_S1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_C1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_S0 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_B1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_D1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_S0 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A2 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_X (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A3 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_C_N (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_SCE (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_C1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_D_N (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_X (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A3 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_A2 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_B (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S0 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A3 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S0 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_B (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A3 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_SCD (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_C (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_C (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_X (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_C1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_S1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_SCD (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_C1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout3_A (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_X (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_X (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A3 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A2 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_X (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_A2 (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_S1 (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_S0 (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_S1 (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_A3 (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_X (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A2 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_X (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A3 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A2 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_B (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_D1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_D_N (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_X (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A2 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A3 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_B (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_X (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_C1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_C (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_C (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_C (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_C1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_C_N (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A0 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A2 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_X (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_D1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout4_A (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone37_C_N (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_X (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_X (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_C_N (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A3 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_C (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A3 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_B (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A3 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_C (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_X (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A3 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_D1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_D_N (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_C (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_S0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_X (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A0 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_C_N (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_S0 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A0 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_C1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_C_N (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_X (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_D1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_D1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_C (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_C1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_C (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_X (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A3 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A3 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_S0 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_C_N (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_B (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_B (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_C1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_X (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_C_N (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_C (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A3 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_S1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_D1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_D1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_D_N (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_S0 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_X (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A2 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_D_N (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_C1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_C (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_SET_B (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_C (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_S1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_X (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_D_N (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_D1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_D1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_A (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_X (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A3 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_S1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_S1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_X (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_D1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_C1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_S0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_S0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_S1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_X (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S0 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A3 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_S1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_X (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_S1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_D1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_D1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_S1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_S1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A3 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_S1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A3 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_X (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_S0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_S1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_S1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_S1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_S1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_D1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_D1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_X (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_B1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A2 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A2 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A2 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_B1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_X (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A2 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_S0 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A0 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_SCD (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_B1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_C_N (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A3 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_S1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_S0 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_S1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_X (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_S0 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_X (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A3 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A2 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S1 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S1 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_S0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_D_N (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_X (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A3 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_S1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_S1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_D1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_S1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_X (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A0 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A3 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_X (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_C_N (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_S0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_D1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_B1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_X (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A3 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_B (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_A (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A3 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_C_N (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_X (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_D1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_SET_B (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_S1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_S0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_C_N (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_X (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A0 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_X (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_S1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_C1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_S0 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S0 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_C (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_X (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_A (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_S1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_A2 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A2 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_S1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_S0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_C1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_B (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_X (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_C (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_B1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_B (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_X (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A3 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_A0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_C (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_A (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_C1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_C (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_B1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone30_C (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_X (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_C (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_C (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_C_N (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_C (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_C1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_D_N (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_X (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_S0 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_S1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A3 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_D1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_C (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone45_A (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_X (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_C (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_S0 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_B1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_C (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_X (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_C1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A3 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S0 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A3 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A2 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_D1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A2 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A3 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_X (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A0 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A3 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A2 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A2 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_X (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A3 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A3 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_X (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A3 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A2 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_A3 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A3 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A2 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A3 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S0 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_D1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_C (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_B (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_X (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A0 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A2 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A3 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A2 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_SCE (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_D1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A2 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_B (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_B (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_B (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_X (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_SCD (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_D_N (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_A1 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A1 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A1 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A2 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_C_N (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_C1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_X (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_S0 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A3 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A2 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_S0 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A0 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_S0 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A2 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_X (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A3 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A3 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_S0 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A2 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A2 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_X (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A3 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S1 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A2 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_S1 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_C1 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A3 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_X (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_D1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A3 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_D1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_X (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S1 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A1 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_S0 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A3 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A1 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_C (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_X (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_S1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_B (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S0 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_C (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_S0 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A2 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_X (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S0 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_X (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A0 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A2 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_C1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A3 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A2 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_C1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_X (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_D1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_C (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A3 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_C (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_D_N (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_C (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_A (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_X (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A0 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A3 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A2 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_S0 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_C (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A3 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_X (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_S1 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A3 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A2 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A0 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A2 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A2 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_S0 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A3 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_A (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_X (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_C_N (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A2 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A2 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_C1 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_B (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_B (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_C1 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge888_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s905_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge848_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_SLEEP_B (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_SLEEP_B (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s922_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s945_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s961_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge854_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge875_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge886_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_SLEEP_B (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_GATE (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge877_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s958_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s959_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s960_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_X (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(clknet_1_0__leaf_net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A2 (.DIODE(clknet_1_0__leaf_net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net604_X (.DIODE(clknet_1_0__leaf_net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_S0 (.DIODE(clknet_1_0__leaf_net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0 (.DIODE(clknet_1_0__leaf_net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S1 (.DIODE(clknet_1_0__leaf_net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net805_X (.DIODE(clknet_1_0__leaf_net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_S0 (.DIODE(clknet_1_1__leaf_net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(clknet_1_1__leaf_net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A0 (.DIODE(clknet_1_1__leaf_net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(clknet_1_1__leaf_net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net380_X (.DIODE(clknet_1_1__leaf_net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A3 (.DIODE(clknet_1_0__leaf_net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S0 (.DIODE(clknet_1_0__leaf_net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_S0 (.DIODE(clknet_1_0__leaf_net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A0 (.DIODE(clknet_1_0__leaf_net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net479_X (.DIODE(clknet_1_0__leaf_net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S1 (.DIODE(clknet_1_1__leaf_net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(clknet_1_1__leaf_net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net951_X (.DIODE(clknet_1_1__leaf_net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net269_A (.DIODE(clknet_0_net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net269_A (.DIODE(clknet_0_net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net269_X (.DIODE(clknet_0_net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A1 (.DIODE(clknet_1_0__leaf_net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A3 (.DIODE(clknet_1_0__leaf_net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_B1 (.DIODE(clknet_1_0__leaf_net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A1 (.DIODE(clknet_1_0__leaf_net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A3 (.DIODE(clknet_1_0__leaf_net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S0 (.DIODE(clknet_1_0__leaf_net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net269_X (.DIODE(clknet_1_0__leaf_net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(clknet_1_0__leaf_net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S1 (.DIODE(clknet_1_0__leaf_net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S0 (.DIODE(clknet_1_0__leaf_net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S0 (.DIODE(clknet_1_0__leaf_net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S0 (.DIODE(clknet_1_0__leaf_net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net767_X (.DIODE(clknet_1_0__leaf_net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_SCE (.DIODE(clknet_1_1__leaf_net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_D1 (.DIODE(clknet_1_1__leaf_net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A3 (.DIODE(clknet_1_1__leaf_net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_S1 (.DIODE(clknet_1_1__leaf_net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_D1 (.DIODE(clknet_1_1__leaf_net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net767_X (.DIODE(clknet_1_1__leaf_net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_B1 (.DIODE(clknet_1_0__leaf_net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A0 (.DIODE(clknet_1_0__leaf_net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A0 (.DIODE(clknet_1_0__leaf_net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(clknet_1_0__leaf_net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(clknet_1_0__leaf_net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net913_X (.DIODE(clknet_1_0__leaf_net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_S0 (.DIODE(clknet_1_1__leaf_net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_D1 (.DIODE(clknet_1_1__leaf_net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A3 (.DIODE(clknet_1_1__leaf_net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S0 (.DIODE(clknet_1_1__leaf_net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(clknet_1_1__leaf_net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S0 (.DIODE(clknet_1_1__leaf_net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A1 (.DIODE(clknet_1_1__leaf_net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net913_X (.DIODE(clknet_1_1__leaf_net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A2 (.DIODE(clknet_1_0__leaf_net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_S0 (.DIODE(clknet_1_0__leaf_net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A3 (.DIODE(clknet_1_0__leaf_net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net706_X (.DIODE(clknet_1_0__leaf_net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A3 (.DIODE(clknet_1_1__leaf_net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S1 (.DIODE(clknet_1_1__leaf_net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_S0 (.DIODE(clknet_1_1__leaf_net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net706_X (.DIODE(clknet_1_1__leaf_net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_B1 (.DIODE(clknet_1_0__leaf_net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A2 (.DIODE(clknet_1_0__leaf_net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_B1 (.DIODE(clknet_1_0__leaf_net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A2 (.DIODE(clknet_1_0__leaf_net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_B1 (.DIODE(clknet_1_0__leaf_net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A3 (.DIODE(clknet_1_0__leaf_net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A2 (.DIODE(clknet_1_0__leaf_net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net343_X (.DIODE(clknet_1_0__leaf_net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A1 (.DIODE(clknet_1_1__leaf_net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A3 (.DIODE(clknet_1_1__leaf_net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A1 (.DIODE(clknet_1_1__leaf_net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A2 (.DIODE(clknet_1_1__leaf_net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A1 (.DIODE(clknet_1_1__leaf_net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A0 (.DIODE(clknet_1_1__leaf_net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S0 (.DIODE(clknet_1_1__leaf_net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net343_X (.DIODE(clknet_1_1__leaf_net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A2 (.DIODE(clknet_1_1__leaf_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A2 (.DIODE(clknet_1_1__leaf_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A3 (.DIODE(clknet_1_1__leaf_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A1 (.DIODE(clknet_1_1__leaf_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A3 (.DIODE(clknet_1_1__leaf_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net354_X (.DIODE(clknet_1_1__leaf_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A1 (.DIODE(clknet_1_0__leaf_net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A2 (.DIODE(clknet_1_0__leaf_net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A1 (.DIODE(clknet_1_0__leaf_net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A0 (.DIODE(clknet_1_0__leaf_net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net232_X (.DIODE(clknet_1_0__leaf_net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A1 (.DIODE(clknet_1_1__leaf_net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_S0 (.DIODE(clknet_1_1__leaf_net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A0 (.DIODE(clknet_1_1__leaf_net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S0 (.DIODE(clknet_1_1__leaf_net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S0 (.DIODE(clknet_1_1__leaf_net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(clknet_1_1__leaf_net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net232_X (.DIODE(clknet_1_1__leaf_net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A2 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A3 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_S0 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer4_X (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A0 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer29_A (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer28_X (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A3 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_S0 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer28_A (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_C1 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone30_X (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_C1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_S0 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_S0 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A3 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A3 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone31_X (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer36_A (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A2 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone37_X (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A1 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A2 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A3 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A3 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A2 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone38_X (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_C1 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A2 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_D1 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A2 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_S0 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone43_X (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_C (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_D1 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A0 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A3 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A3 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone44_X (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_B1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_C (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_SCE (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone45_X (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout2_X (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_D_N (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_B1 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_C1 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A1 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A0 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_C1 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A2 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S0 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_B1 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout3_X (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A2 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A3 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A3 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A2 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_S1 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone37_A (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A2 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout4_X (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_C_N (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_S0 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_C1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S0 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_B (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_S1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_D1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_C (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_C (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout5_X (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A3 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A2 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone30_B (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_B (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_A (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A2 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_D1 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_D1 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_D1 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_B1 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net78));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net86),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(net1110),
    .X(net1109));
 sky130_fd_sc_hd__mux4_1 clone32 (.A0(net989),
    .A1(net83),
    .A2(net85),
    .A3(net1001),
    .S0(net69),
    .S1(net1013),
    .X(net1110));
 sky130_fd_sc_hd__mux4_1 clone33 (.A0(net992),
    .A1(net75),
    .A2(net80),
    .A3(net73),
    .S0(net74),
    .S1(net1002),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer37 (.A(net69),
    .X(net1112));
 sky130_fd_sc_hd__and3_1 clone39 (.A(net1013),
    .B(net1040),
    .C(net1023),
    .X(net1113));
 sky130_fd_sc_hd__and3_1 clone40 (.A(net1040),
    .B(net1038),
    .C(net1027),
    .X(net1114));
 sky130_fd_sc_hd__or4bb_1 clone42 (.A(net1105),
    .B(net85),
    .C_N(net1106),
    .D_N(net1104),
    .X(net1115));
 sky130_fd_sc_hd__a2111o_1 clone46 (.A1(net103),
    .A2(net862),
    .B1(net871),
    .C1(net1103),
    .D1(net101),
    .X(net1116));
 sky130_fd_sc_hd__mux4_1 clone47 (.A0(net11),
    .A1(net21),
    .A2(net1128),
    .A3(net22),
    .S0(net14),
    .S1(net12),
    .X(net1117));
 sky130_fd_sc_hd__mux4_1 clone48 (.A0(net898),
    .A1(net899),
    .A2(net3),
    .A3(net897),
    .S0(net0),
    .S1(net890),
    .X(net1118));
 sky130_fd_sc_hd__and3_1 clone49 (.A(net1106),
    .B(net1046),
    .C(net73),
    .X(net1119));
 sky130_fd_sc_hd__mux4_1 clone50 (.A0(net991),
    .A1(net18),
    .A2(net1107),
    .A3(net23),
    .S0(net887),
    .S1(net987),
    .X(net1120));
 sky130_fd_sc_hd__mux4_1 clone51 (.A0(net11),
    .A1(net21),
    .A2(net1128),
    .A3(net22),
    .S0(net14),
    .S1(net12),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer52 (.A(net73),
    .X(net1122));
 sky130_fd_sc_hd__and3_1 clone53 (.A(net1124),
    .B(net1027),
    .C(net1040),
    .X(net1123));
 sky130_fd_sc_hd__and3_1 clone54 (.A(net1013),
    .B(net1040),
    .C(net1023),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer55 (.A(net24),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer56 (.A(net46),
    .X(net1126));
 sky130_fd_sc_hd__mux4_1 clone57 (.A0(net45),
    .A1(net1085),
    .A2(net939),
    .A3(net27),
    .S0(net30),
    .S1(net44),
    .X(net1127));
 sky130_fd_sc_hd__a2111o_1 clone58 (.A1(net17),
    .A2(net11),
    .B1(net10),
    .C1(net1042),
    .D1(net1107),
    .X(net1128));
 sky130_fd_sc_hd__and3_1 clone59 (.A(net997),
    .B(net1013),
    .C(net1043),
    .X(net1129));
 sky130_fd_sc_hd__mux4_1 clone60 (.A0(net991),
    .A1(net18),
    .A2(net1107),
    .A3(net23),
    .S0(net887),
    .S1(net987),
    .X(net1130));
 sky130_fd_sc_hd__clkbuf_1 clone61 (.A(net24),
    .X(net1131));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
