module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net165;
 wire net176;
 wire net703;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net818;
 wire clknet_1_0__leaf_net818;
 wire clknet_1_1__leaf_net818;
 wire clknet_0_net615;
 wire clknet_1_0__leaf_net615;
 wire clknet_1_1__leaf_net615;
 wire clknet_0_net817;
 wire clknet_1_0__leaf_net817;
 wire clknet_1_1__leaf_net817;
 wire clknet_0_net608;
 wire clknet_1_0__leaf_net608;
 wire clknet_1_1__leaf_net608;
 wire clknet_0_net600;
 wire clknet_1_0__leaf_net600;
 wire clknet_1_1__leaf_net600;
 wire clknet_0_net711;
 wire clknet_1_0__leaf_net711;
 wire clknet_1_1__leaf_net711;
 wire clknet_0_net611;
 wire clknet_1_0__leaf_net611;
 wire clknet_1_1__leaf_net611;
 wire clknet_0_net577;
 wire clknet_1_0__leaf_net577;
 wire clknet_1_1__leaf_net577;
 wire clknet_0_net798;
 wire clknet_1_0__leaf_net798;
 wire clknet_1_1__leaf_net798;
 wire clknet_0_net511;
 wire clknet_1_0__leaf_net511;
 wire clknet_1_1__leaf_net511;
 wire clknet_0_net797;
 wire clknet_1_0__leaf_net797;
 wire clknet_1_1__leaf_net797;
 wire clknet_0_net602;
 wire clknet_1_0__leaf_net602;
 wire clknet_1_1__leaf_net602;
 wire clknet_0_net495;
 wire clknet_1_0__leaf_net495;
 wire clknet_1_1__leaf_net495;
 wire clknet_0_net502;
 wire clknet_1_0__leaf_net502;
 wire clknet_1_1__leaf_net502;
 wire clknet_0_net796;
 wire clknet_1_0__leaf_net796;
 wire clknet_1_1__leaf_net796;
 wire clknet_0_net777;
 wire clknet_1_0__leaf_net777;
 wire clknet_1_1__leaf_net777;
 wire clknet_0_net398;
 wire clknet_1_0__leaf_net398;
 wire clknet_1_1__leaf_net398;
 wire clknet_0_net610;
 wire clknet_1_0__leaf_net610;
 wire clknet_1_1__leaf_net610;
 wire clknet_0_net420;
 wire clknet_1_0__leaf_net420;
 wire clknet_1_1__leaf_net420;
 wire clknet_0_net391;
 wire clknet_1_0__leaf_net391;
 wire clknet_1_1__leaf_net391;
 wire clknet_0_net389;
 wire clknet_1_0__leaf_net389;
 wire clknet_1_1__leaf_net389;
 wire clknet_0_net776;
 wire clknet_1_0__leaf_net776;
 wire clknet_1_1__leaf_net776;
 wire clknet_0_net775;
 wire clknet_1_0__leaf_net775;
 wire clknet_1_1__leaf_net775;
 wire clknet_0_net595;
 wire clknet_1_0__leaf_net595;
 wire clknet_1_1__leaf_net595;
 wire clknet_0_net901;
 wire clknet_1_0__leaf_net901;
 wire clknet_1_1__leaf_net901;
 wire clknet_0_net186;
 wire clknet_1_0__leaf_net186;
 wire clknet_1_1__leaf_net186;
 wire clknet_0_net910;
 wire clknet_1_0__leaf_net910;
 wire clknet_1_1__leaf_net910;
 wire clknet_0_net179;
 wire clknet_1_0__leaf_net179;
 wire clknet_1_1__leaf_net179;
 wire clknet_0_net180;
 wire clknet_1_0__leaf_net180;
 wire clknet_1_1__leaf_net180;
 wire clknet_0_net759;
 wire clknet_1_0__leaf_net759;
 wire clknet_1_1__leaf_net759;
 wire clknet_0_net924;
 wire clknet_1_0__leaf_net924;
 wire clknet_1_1__leaf_net924;
 wire clknet_0_net905;
 wire clknet_1_0__leaf_net905;
 wire clknet_1_1__leaf_net905;
 wire clknet_0_net177;
 wire clknet_1_0__leaf_net177;
 wire clknet_1_1__leaf_net177;
 wire clknet_0_net902;
 wire clknet_1_0__leaf_net902;
 wire clknet_1_1__leaf_net902;
 wire clknet_0_net709;
 wire clknet_1_0__leaf_net709;
 wire clknet_1_1__leaf_net709;
 wire clknet_0_net758;
 wire clknet_1_0__leaf_net758;
 wire clknet_1_1__leaf_net758;
 wire clknet_0_net281;
 wire clknet_1_0__leaf_net281;
 wire clknet_1_1__leaf_net281;
 wire clknet_0_net911;
 wire clknet_1_0__leaf_net911;
 wire clknet_1_1__leaf_net911;
 wire clknet_0_net276;
 wire clknet_1_0__leaf_net276;
 wire clknet_1_1__leaf_net276;
 wire clknet_0_net170;
 wire clknet_1_0__leaf_net170;
 wire clknet_1_1__leaf_net170;
 wire clknet_0_net744;
 wire clknet_1_0__leaf_net744;
 wire clknet_1_1__leaf_net744;
 wire clknet_0_net532;
 wire clknet_1_0__leaf_net532;
 wire clknet_1_1__leaf_net532;
 wire clknet_0_net879;
 wire clknet_1_0__leaf_net879;
 wire clknet_1_1__leaf_net879;
 wire clknet_0_net710;
 wire clknet_1_0__leaf_net710;
 wire clknet_1_1__leaf_net710;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;

 sky130_fd_sc_hd__a21bo_2 c100 (.A1(net1002),
    .A2(net11),
    .B1_N(net1000),
    .X(net37));
 sky130_fd_sc_hd__a41o_1 c101 (.A1(net36),
    .A2(net35),
    .A3(net11),
    .A4(net834),
    .B1(net34),
    .X(net38));
 sky130_fd_sc_hd__a21bo_1 c102 (.A1(net37),
    .A2(net30),
    .B1_N(net29),
    .X(net39));
 sky130_fd_sc_hd__a31o_1 c103 (.A1(net34),
    .A2(net32),
    .A3(net35),
    .B1(net972),
    .X(net40));
 sky130_fd_sc_hd__mux4_2 c104 (.A0(net38),
    .A1(net33),
    .A2(net1019),
    .A3(net24),
    .S0(net837),
    .S1(net35),
    .X(net41));
 sky130_fd_sc_hd__a41o_4 c105 (.A1(net41),
    .A2(net29),
    .A3(net31),
    .A4(net36),
    .B1(net1004),
    .X(net42));
 sky130_fd_sc_hd__mux4_2 c106 (.A0(net31),
    .A1(net38),
    .A2(net42),
    .A3(net8),
    .S0(net951),
    .S1(net1034),
    .X(net43));
 sky130_fd_sc_hd__a41o_4 c107 (.A1(net28),
    .A2(net871),
    .A3(net42),
    .A4(net856),
    .B1(net43),
    .X(net884));
 sky130_fd_sc_hd__mux4_2 c108 (.A0(net11),
    .A1(net34),
    .A2(net41),
    .A3(net33),
    .S0(net951),
    .S1(net972),
    .X(net44));
 sky130_fd_sc_hd__a41o_1 c109 (.A1(net41),
    .A2(net38),
    .A3(net44),
    .A4(net7),
    .B1(net43),
    .X(net45));
 sky130_fd_sc_hd__mux4_1 c110 (.A0(net997),
    .A1(net871),
    .A2(net31),
    .A3(net35),
    .S0(net971),
    .S1(net1018),
    .X(net46));
 sky130_fd_sc_hd__a21bo_1 c111 (.A1(net862),
    .A2(net6),
    .B1_N(net1007),
    .X(net47));
 sky130_fd_sc_hd__a31o_1 c112 (.A1(net37),
    .A2(net6),
    .A3(net860),
    .B1(net865),
    .X(net48));
 sky130_fd_sc_hd__a21bo_2 c113 (.A1(net844),
    .A2(net862),
    .B1_N(net1021),
    .X(net49));
 sky130_fd_sc_hd__a21bo_1 c114 (.A1(net20),
    .A2(net9),
    .B1_N(net37),
    .X(net50));
 sky130_fd_sc_hd__a31o_1 c115 (.A1(net48),
    .A2(net46),
    .A3(net865),
    .B1(net44),
    .X(net51));
 sky130_fd_sc_hd__a31o_1 c116 (.A1(net990),
    .A2(net25),
    .A3(net50),
    .B1(net1013),
    .X(net52));
 sky130_fd_sc_hd__a21bo_1 c117 (.A1(net51),
    .A2(net48),
    .B1_N(net18),
    .X(net53));
 sky130_fd_sc_hd__a21bo_2 c118 (.A1(net6),
    .A2(net50),
    .B1_N(net1018),
    .X(net894));
 sky130_fd_sc_hd__a41o_1 c119 (.A1(net9),
    .A2(net49),
    .A3(net954),
    .A4(net971),
    .B1(net1015),
    .X(net54));
 sky130_fd_sc_hd__a41o_1 c120 (.A1(net1007),
    .A2(net51),
    .A3(net18),
    .A4(net971),
    .B1(net865),
    .X(net55));
 sky130_fd_sc_hd__a41o_1 c121 (.A1(net18),
    .A2(net25),
    .A3(net55),
    .A4(net51),
    .B1(net954),
    .X(net913));
 sky130_fd_sc_hd__a21bo_1 c122 (.A1(net833),
    .A2(net913),
    .B1_N(net49),
    .X(net56));
 sky130_fd_sc_hd__mux4_1 c123 (.A0(net56),
    .A1(net54),
    .A2(net1018),
    .A3(net51),
    .S0(net833),
    .S1(net1044),
    .X(net57));
 sky130_fd_sc_hd__a21bo_1 c124 (.A1(net31),
    .A2(net47),
    .B1_N(net954),
    .X(net58));
 sky130_fd_sc_hd__a41o_1 c125 (.A1(net1015),
    .A2(net55),
    .A3(net47),
    .A4(net954),
    .B1(net58),
    .X(net59));
 sky130_fd_sc_hd__mux4_2 c126 (.A0(net55),
    .A1(net52),
    .A2(net954),
    .A3(net6),
    .S0(net1021),
    .S1(net751),
    .X(net60));
 sky130_fd_sc_hd__mux4_2 c127 (.A0(net871),
    .A1(net51),
    .A2(net60),
    .A3(net9),
    .S0(net1006),
    .S1(net954),
    .X(net61));
 sky130_fd_sc_hd__a41o_1 c128 (.A1(net60),
    .A2(net48),
    .A3(net954),
    .A4(net59),
    .B1(net1044),
    .X(net62));
 sky130_fd_sc_hd__mux4_1 c129 (.A0(net44),
    .A1(net60),
    .A2(net62),
    .A3(net972),
    .S0(net49),
    .S1(net61),
    .X(net63));
 sky130_fd_sc_hd__mux4_1 c130 (.A0(net46),
    .A1(net62),
    .A2(net56),
    .A3(net50),
    .S0(net6),
    .S1(net927),
    .X(net64));
 sky130_fd_sc_hd__sdfbbn_1 c131 (.CLK_N(clknet_4_4_0_clk),
    .D(net60),
    .RESET_B(net61),
    .SCD(net46),
    .SCE(net9),
    .SET_B(net927),
    .Q(net66),
    .Q_N(net65));
 sky130_fd_sc_hd__a21bo_2 c132 (.A1(net1019),
    .A2(net1016),
    .B1_N(net995),
    .X(net67));
 sky130_fd_sc_hd__a31o_4 c133 (.A1(net67),
    .A2(net703),
    .A3(net1002),
    .B1(net1023),
    .X(net68));
 sky130_fd_sc_hd__a21bo_2 c134 (.A1(net1018),
    .A2(net996),
    .B1_N(net1022),
    .X(net69));
 sky130_fd_sc_hd__a21bo_1 c135 (.A1(net1002),
    .A2(net1005),
    .B1_N(net995),
    .X(net70));
 sky130_fd_sc_hd__a21bo_2 c136 (.A1(net1002),
    .A2(net1016),
    .B1_N(net998),
    .X(net71));
 sky130_fd_sc_hd__a21bo_2 c137 (.A1(net995),
    .A2(net996),
    .B1_N(net991),
    .X(net72));
 sky130_fd_sc_hd__a21bo_2 c138 (.A1(net1014),
    .A2(net1021),
    .B1_N(net67),
    .X(net73));
 sky130_fd_sc_hd__a21bo_4 c139 (.A1(net67),
    .A2(net995),
    .B1_N(net991),
    .X(net74));
 sky130_fd_sc_hd__a21bo_2 c140 (.A1(net1025),
    .A2(net703),
    .B1_N(net984),
    .X(net75));
 sky130_fd_sc_hd__a41o_4 c141 (.A1(net983),
    .A2(net995),
    .A3(net1016),
    .A4(net75),
    .B1(net998),
    .X(net76));
 sky130_fd_sc_hd__a41o_1 c142 (.A1(net1023),
    .A2(net1024),
    .A3(net1002),
    .A4(net983),
    .B1(net991),
    .X(net77));
 sky130_fd_sc_hd__xnor2_4 c143 (.A(net1012),
    .B(net1025),
    .Y(net78));
 sky130_fd_sc_hd__a21bo_4 c144 (.A1(net76),
    .A2(net1009),
    .B1_N(net78),
    .X(net79));
 sky130_fd_sc_hd__a21bo_4 c145 (.A1(net993),
    .A2(net67),
    .B1_N(net1004),
    .X(net80));
 sky130_fd_sc_hd__a21bo_4 c146 (.A1(net80),
    .A2(net1024),
    .B1_N(net980),
    .X(net81));
 sky130_fd_sc_hd__mux4_2 c147 (.A0(net991),
    .A1(net1002),
    .A2(net79),
    .A3(net81),
    .S0(net998),
    .S1(net983),
    .X(net82));
 sky130_fd_sc_hd__a21bo_1 c148 (.A1(net993),
    .A2(net969),
    .B1_N(net980),
    .X(net83));
 sky130_fd_sc_hd__mux4_2 c149 (.A0(net80),
    .A1(net1024),
    .A2(net827),
    .A3(net1003),
    .S0(net1005),
    .S1(net71),
    .X(net84));
 sky130_fd_sc_hd__mux4_2 c150 (.A0(net71),
    .A1(net1012),
    .A2(net84),
    .A3(net1009),
    .S0(net980),
    .S1(net74),
    .X(net85));
 sky130_fd_sc_hd__a21bo_2 c151 (.A1(net84),
    .A2(net85),
    .B1_N(net67),
    .X(net86));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net85),
    .A1(net83),
    .A2(net983),
    .A3(net84),
    .S0(net79),
    .S1(net86),
    .X(net87));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net87),
    .A1(net84),
    .A2(net85),
    .A3(net86),
    .S0(net994),
    .S1(net1024),
    .X(net88));
 sky130_fd_sc_hd__a41o_1 c154 (.A1(net847),
    .A2(net78),
    .A3(net1005),
    .A4(net1013),
    .B1(net995),
    .X(net903));
 sky130_fd_sc_hd__a21bo_1 c155 (.A1(net998),
    .A2(net86),
    .B1_N(net68),
    .X(net89));
 sky130_fd_sc_hd__a21bo_1 c156 (.A1(net854),
    .A2(net1015),
    .B1_N(net84),
    .X(net90));
 sky130_fd_sc_hd__a31o_4 c157 (.A1(net1019),
    .A2(net83),
    .A3(net1013),
    .B1(net853),
    .X(net91));
 sky130_fd_sc_hd__a31o_1 c158 (.A1(net834),
    .A2(net838),
    .A3(net1010),
    .B1(net981),
    .X(net92));
 sky130_fd_sc_hd__a41o_1 c159 (.A1(net90),
    .A2(net836),
    .A3(net827),
    .A4(net969),
    .B1(net1016),
    .X(net93));
 sky130_fd_sc_hd__a21bo_1 c160 (.A1(net838),
    .A2(net91),
    .B1_N(net93),
    .X(net94));
 sky130_fd_sc_hd__a21bo_2 c161 (.A1(net93),
    .A2(net836),
    .B1_N(net81),
    .X(net95));
 sky130_fd_sc_hd__mux4_2 c162 (.A0(net95),
    .A1(net92),
    .A2(net1014),
    .A3(net837),
    .S0(net981),
    .S1(net998),
    .X(net96));
 sky130_fd_sc_hd__a41o_2 c163 (.A1(net89),
    .A2(net983),
    .A3(net91),
    .A4(net838),
    .B1(net981),
    .X(net881));
 sky130_fd_sc_hd__a41o_2 c164 (.A1(net703),
    .A2(net853),
    .A3(net1010),
    .A4(net1003),
    .B1(net95),
    .X(net97));
 sky130_fd_sc_hd__a41o_4 c165 (.A1(net969),
    .A2(net97),
    .A3(net836),
    .A4(net844),
    .B1(net982),
    .X(net98));
 sky130_fd_sc_hd__a41o_1 c166 (.A1(net96),
    .A2(net1025),
    .A3(net98),
    .A4(net837),
    .B1(net833),
    .X(net99));
 sky130_fd_sc_hd__a41o_2 c167 (.A1(net99),
    .A2(net94),
    .A3(net84),
    .A4(net96),
    .B1(net98),
    .X(net100));
 sky130_fd_sc_hd__a41o_2 c168 (.A1(net89),
    .A2(net100),
    .A3(net92),
    .A4(net1018),
    .B1(net960),
    .X(net101));
 sky130_fd_sc_hd__mux4_2 c169 (.A0(net96),
    .A1(net99),
    .A2(net91),
    .A3(net100),
    .S0(net97),
    .S1(net847),
    .X(net102));
 sky130_fd_sc_hd__a41o_4 c170 (.A1(net94),
    .A2(net89),
    .A3(net100),
    .A4(net1019),
    .B1(net97),
    .X(net103));
 sky130_fd_sc_hd__a41o_2 c171 (.A1(net846),
    .A2(net90),
    .A3(net960),
    .A4(net949),
    .B1(net1004),
    .X(net104));
 sky130_fd_sc_hd__mux4_2 c172 (.A0(net102),
    .A1(net100),
    .A2(net827),
    .A3(net104),
    .S0(net97),
    .S1(net949),
    .X(net919));
 sky130_fd_sc_hd__mux4_2 c173 (.A0(net104),
    .A1(net95),
    .A2(net943),
    .A3(net847),
    .S0(net949),
    .S1(net100),
    .X(net105));
 sky130_fd_sc_hd__mux4_2 c174 (.A0(net100),
    .A1(net980),
    .A2(net949),
    .A3(net991),
    .S0(net84),
    .S1(net936),
    .X(net106));
 sky130_fd_sc_hd__mux4_2 c175 (.A0(net936),
    .A1(net841),
    .A2(net106),
    .A3(net943),
    .S0(net961),
    .S1(net104),
    .X(net107));
 sky130_fd_sc_hd__a41o_1 c176 (.A1(net827),
    .A2(net104),
    .A3(net856),
    .A4(net990),
    .B1(net1023),
    .X(net108));
 sky130_fd_sc_hd__a21bo_1 c177 (.A1(net94),
    .A2(net1),
    .B1_N(net1004),
    .X(net914));
 sky130_fd_sc_hd__a21bo_2 c178 (.A1(net83),
    .A2(net870),
    .B1_N(net86),
    .X(net109));
 sky130_fd_sc_hd__a41o_2 c179 (.A1(net869),
    .A2(net106),
    .A3(net991),
    .A4(net847),
    .B1(net1000),
    .X(net110));
 sky130_fd_sc_hd__a21bo_2 c180 (.A1(net952),
    .A2(net2),
    .B1_N(net1010),
    .X(net111));
 sky130_fd_sc_hd__a41o_1 c181 (.A1(net1003),
    .A2(net840),
    .A3(net856),
    .A4(net873),
    .B1(net943),
    .X(net112));
 sky130_fd_sc_hd__a21bo_4 c182 (.A1(net844),
    .A2(net1),
    .B1_N(net1012),
    .X(net113));
 sky130_fd_sc_hd__a21bo_1 c183 (.A1(net97),
    .A2(net858),
    .B1_N(net109),
    .X(net114));
 sky130_fd_sc_hd__a41o_1 c184 (.A1(net114),
    .A2(net81),
    .A3(net110),
    .A4(net852),
    .B1(net847),
    .X(net115));
 sky130_fd_sc_hd__a31o_4 c185 (.A1(net113),
    .A2(net846),
    .A3(net1002),
    .B1(net114),
    .X(net116));
 sky130_fd_sc_hd__a21bo_1 c186 (.A1(net79),
    .A2(net107),
    .B1_N(net114),
    .X(net117));
 sky130_fd_sc_hd__a41o_1 c187 (.A1(net849),
    .A2(net870),
    .A3(net113),
    .A4(net116),
    .B1(net995),
    .X(net118));
 sky130_fd_sc_hd__a21bo_1 c188 (.A1(net112),
    .A2(net949),
    .B1_N(net991),
    .X(net119));
 sky130_fd_sc_hd__a21bo_2 c189 (.A1(net84),
    .A2(net2),
    .B1_N(net953),
    .X(net120));
 sky130_fd_sc_hd__a21bo_2 c190 (.A1(net120),
    .A2(net114),
    .B1_N(net119),
    .X(net121));
 sky130_fd_sc_hd__a41o_2 c191 (.A1(net119),
    .A2(net120),
    .A3(net865),
    .A4(net1010),
    .B1(net1007),
    .X(net122));
 sky130_fd_sc_hd__a41o_2 c192 (.A1(net116),
    .A2(net114),
    .A3(net935),
    .A4(net1015),
    .B1(net953),
    .X(net123));
 sky130_fd_sc_hd__a41o_1 c193 (.A1(net935),
    .A2(net117),
    .A3(net119),
    .A4(net121),
    .B1(net108),
    .X(net124));
 sky130_fd_sc_hd__a41o_2 c194 (.A1(net118),
    .A2(net115),
    .A3(net120),
    .A4(net124),
    .B1(net1007),
    .X(net909));
 sky130_fd_sc_hd__a21bo_2 c195 (.A1(net111),
    .A2(net121),
    .B1_N(net935),
    .X(net125));
 sky130_fd_sc_hd__mux4_2 c196 (.A0(net124),
    .A1(net119),
    .A2(net123),
    .A3(net863),
    .S0(net120),
    .S1(net125),
    .X(net126));
 sky130_fd_sc_hd__mux4_2 c197 (.A0(net93),
    .A1(net108),
    .A2(net97),
    .A3(net111),
    .S0(net113),
    .S1(net116),
    .X(net127));
 sky130_fd_sc_hd__a21bo_1 c198 (.A1(net111),
    .A2(net74),
    .B1_N(net109),
    .X(net128));
 sky130_fd_sc_hd__a21bo_4 c199 (.A1(net21),
    .A2(net79),
    .B1_N(net109),
    .X(net891));
 sky130_fd_sc_hd__a21bo_4 c200 (.A1(net874),
    .A2(net868),
    .B1_N(net1007),
    .X(net129));
 sky130_fd_sc_hd__a21bo_1 c201 (.A1(net5),
    .A2(net129),
    .B1_N(net992),
    .X(net130));
 sky130_fd_sc_hd__a41o_1 c202 (.A1(net949),
    .A2(net128),
    .A3(net14),
    .A4(net104),
    .B1(net1030),
    .X(net131));
 sky130_fd_sc_hd__a41o_1 c203 (.A1(net106),
    .A2(net124),
    .A3(net1039),
    .A4(net130),
    .B1(net849),
    .X(net132));
 sky130_fd_sc_hd__a41o_1 c204 (.A1(net103),
    .A2(net833),
    .A3(net129),
    .A4(net1045),
    .B1(net1000),
    .X(net133));
 sky130_fd_sc_hd__a21bo_2 c205 (.A1(net845),
    .A2(net115),
    .B1_N(net0),
    .X(net134));
 sky130_fd_sc_hd__a41o_1 c206 (.A1(net74),
    .A2(net134),
    .A3(net842),
    .A4(net1045),
    .B1(net81),
    .X(net135));
 sky130_fd_sc_hd__mux4_1 c207 (.A0(net14),
    .A1(net113),
    .A2(net134),
    .A3(net103),
    .S0(net992),
    .S1(net1039),
    .X(net136));
 sky130_fd_sc_hd__a21bo_1 c208 (.A1(net130),
    .A2(net79),
    .B1_N(net20),
    .X(net137));
 sky130_fd_sc_hd__a21bo_2 c209 (.A1(net129),
    .A2(net863),
    .B1_N(net957),
    .X(net138));
 sky130_fd_sc_hd__sdfbbn_2 c210 (.CLK_N(clknet_4_1_0_clk),
    .D(net134),
    .RESET_B(net874),
    .SCD(net957),
    .SCE(net136),
    .SET_B(net132),
    .Q(net888),
    .Q_N(net139));
 sky130_fd_sc_hd__mux4_2 c211 (.A0(net842),
    .A1(net112),
    .A2(net123),
    .A3(net1010),
    .S0(net1045),
    .S1(net957),
    .X(net140));
 sky130_fd_sc_hd__a41o_1 c212 (.A1(net841),
    .A2(net138),
    .A3(net140),
    .A4(net957),
    .B1(net953),
    .X(net141));
 sky130_fd_sc_hd__mux4_2 c213 (.A0(net133),
    .A1(net20),
    .A2(net5),
    .A3(net14),
    .S0(net24),
    .S1(net140),
    .X(net142));
 sky130_fd_sc_hd__mux4_1 c214 (.A0(net128),
    .A1(net132),
    .A2(net140),
    .A3(net14),
    .S0(net123),
    .S1(net957),
    .X(net143));
 sky130_fd_sc_hd__mux4_1 c215 (.A0(net141),
    .A1(net21),
    .A2(net142),
    .A3(net958),
    .S0(net983),
    .S1(net111),
    .X(net144));
 sky130_fd_sc_hd__a41o_1 c216 (.A1(net140),
    .A2(net837),
    .A3(net957),
    .A4(net1045),
    .B1(net753),
    .X(net145));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(net135),
    .A1(net957),
    .A2(net142),
    .A3(net133),
    .S0(net140),
    .S1(net1049),
    .X(net146));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(net145),
    .A1(net140),
    .A2(net891),
    .A3(net23),
    .S0(net957),
    .S1(net753),
    .X(net147));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net136),
    .A1(net10),
    .A2(net142),
    .A3(net1010),
    .S0(net111),
    .S1(net989),
    .X(net148));
 sky130_fd_sc_hd__a41o_4 c220 (.A1(net140),
    .A2(net1044),
    .A3(net26),
    .A4(net138),
    .B1(net981),
    .X(net880));
 sky130_fd_sc_hd__sdfbbp_1 c221 (.CLK(clknet_4_4_0_clk),
    .D(net141),
    .RESET_B(net1007),
    .SCD(net37),
    .SCE(net1038),
    .SET_B(net32),
    .Q(net898),
    .Q_N(net149));
 sky130_fd_sc_hd__a41o_1 c222 (.A1(net958),
    .A2(net943),
    .A3(net972),
    .A4(net989),
    .B1(net754),
    .X(net150));
 sky130_fd_sc_hd__sdfbbn_1 c223 (.CLK_N(clknet_4_5_0_clk),
    .D(net45),
    .RESET_B(net142),
    .SCD(net109),
    .SCE(net1000),
    .SET_B(net68),
    .Q(net152),
    .Q_N(net151));
 sky130_fd_sc_hd__mux4_1 c224 (.A0(net124),
    .A1(net880),
    .A2(net109),
    .A3(net149),
    .S0(net831),
    .S1(net753),
    .X(net153));
 sky130_fd_sc_hd__a41o_4 c225 (.A1(net884),
    .A2(net951),
    .A3(net664),
    .A4(net754),
    .B1(net755),
    .X(net154));
 sky130_fd_sc_hd__mux4_2 c226 (.A0(net32),
    .A1(net150),
    .A2(net898),
    .A3(net154),
    .S0(net2),
    .S1(net755),
    .X(net155));
 sky130_fd_sc_hd__mux4_1 c227 (.A0(net27),
    .A1(net874),
    .A2(net1015),
    .A3(net997),
    .S0(net664),
    .S1(net755),
    .X(net156));
 sky130_fd_sc_hd__mux4_2 c228 (.A0(net24),
    .A1(net26),
    .A2(net101),
    .A3(net943),
    .S0(net1000),
    .S1(net755),
    .X(net157));
 sky130_fd_sc_hd__mux4_1 c229 (.A0(net43),
    .A1(net150),
    .A2(net16),
    .A3(net101),
    .S0(net1013),
    .S1(net972),
    .X(net158));
 sky130_fd_sc_hd__a41o_1 c230 (.A1(net117),
    .A2(net129),
    .A3(net1033),
    .A4(net45),
    .B1(net151),
    .X(net159));
 sky130_fd_sc_hd__mux4_1 c231 (.A0(net113),
    .A1(net960),
    .A2(net863),
    .A3(net149),
    .S0(net1024),
    .S1(net957),
    .X(net160));
 sky130_fd_sc_hd__a41o_1 c232 (.A1(net156),
    .A2(net40),
    .A3(net26),
    .A4(net1007),
    .B1(net754),
    .X(net161));
 sky130_fd_sc_hd__sdfbbn_2 c233 (.CLK_N(clknet_4_5_0_clk),
    .D(net161),
    .RESET_B(net142),
    .SCD(net116),
    .SCE(net981),
    .SET_B(net754),
    .Q(net904),
    .Q_N(net162));
 sky130_fd_sc_hd__a41o_1 c234 (.A1(net157),
    .A2(net42),
    .A3(net943),
    .A4(net834),
    .B1(net880),
    .X(net163));
 sky130_fd_sc_hd__mux4_1 c235 (.A0(net158),
    .A1(net140),
    .A2(net162),
    .A3(net151),
    .S0(net113),
    .S1(net154),
    .X(net164));
 sky130_fd_sc_hd__mux4_2 c236 (.A0(net155),
    .A1(net149),
    .A2(net162),
    .A3(net156),
    .S0(net664),
    .X(net674));
 sky130_fd_sc_hd__mux4_1 c237 (.A0(net2),
    .A1(net150),
    .A2(net904),
    .A3(net27),
    .S0(net837),
    .S1(net113),
    .X(net166));
 sky130_fd_sc_hd__mux4_1 c238 (.A0(net166),
    .A1(net838),
    .A2(net158),
    .A3(net164),
    .S0(net1011),
    .S1(net162),
    .X(net167));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net164),
    .A1(net113),
    .A2(net166),
    .A3(net1029),
    .S0(net35),
    .S1(net675),
    .X(net168));
 sky130_fd_sc_hd__mux4_1 c240 (.A0(net1033),
    .A1(net904),
    .A2(net161),
    .A3(net880),
    .S0(net117),
    .S1(net675),
    .X(net169));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(net115),
    .A1(net26),
    .A2(net868),
    .A3(net15),
    .S0(net756),
    .S1(clknet_1_0__leaf_net758),
    .X(net170));
 sky130_fd_sc_hd__mux4_2 c242 (.A0(net834),
    .A1(net50),
    .A2(net25),
    .A3(net1015),
    .S0(net674),
    .S1(net751),
    .X(net171));
 sky130_fd_sc_hd__mux4_2 c243 (.A0(net865),
    .A1(net54),
    .A2(net898),
    .A3(net1024),
    .S0(net971),
    .S1(net25),
    .X(net885));
 sky130_fd_sc_hd__mux4_1 c244 (.A0(net854),
    .A1(net160),
    .A2(net139),
    .A3(net31),
    .S0(net931),
    .S1(net1038),
    .X(net172));
 sky130_fd_sc_hd__sdfbbp_1 c245 (.CLK(clknet_4_1_0_clk),
    .D(net913),
    .RESET_B(net931),
    .SCD(net29),
    .SCE(net674),
    .SET_B(clknet_1_0__leaf_net759),
    .Q(net174),
    .Q_N(net173));
 sky130_fd_sc_hd__mux4_1 c246 (.A0(net860),
    .A1(net981),
    .A2(net149),
    .A3(net931),
    .S0(net138),
    .S1(clknet_1_0__leaf_net759),
    .X(net175));
 sky130_fd_sc_hd__mux4_1 c247 (.A0(net61),
    .A1(net171),
    .A2(net1021),
    .A3(net880),
    .S1(clknet_1_1__leaf_net759),
    .X(net709));
 sky130_fd_sc_hd__mux4_1 c248 (.A0(net138),
    .A1(net943),
    .A2(net173),
    .A3(net991),
    .S0(net1023),
    .S1(clknet_1_0__leaf_net759),
    .X(net905));
 sky130_fd_sc_hd__mux4_1 c249 (.A0(net174),
    .A1(net53),
    .A2(net49),
    .A3(net25),
    .S0(net1018),
    .S1(clknet_1_0__leaf_net759),
    .X(net924));
 sky130_fd_sc_hd__mux4_1 c250 (.A0(net29),
    .A1(clknet_1_1__leaf_net905),
    .A2(net171),
    .A3(net52),
    .S0(net898),
    .S1(net112),
    .X(net902));
 sky130_fd_sc_hd__mux4_1 c251 (.A0(net25),
    .A1(net157),
    .A2(net59),
    .A3(clknet_1_0__leaf_net902),
    .S0(clknet_1_1__leaf_net905),
    .S1(clknet_1_0__leaf_net709),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 c252 (.A0(net833),
    .A1(clknet_1_0__leaf_net905),
    .A2(net20),
    .A3(net880),
    .S0(net954),
    .S1(net981),
    .X(net178));
 sky130_fd_sc_hd__mux4_1 c253 (.A0(net54),
    .A1(net885),
    .A2(net20),
    .A3(net1044),
    .S0(net981),
    .S1(clknet_1_0__leaf_net901),
    .X(net179));
 sky130_fd_sc_hd__mux4_1 c254 (.A0(clknet_1_0__leaf_net179),
    .A1(net981),
    .A2(net60),
    .A3(net1015),
    .S0(clknet_1_0__leaf_net709),
    .S1(clknet_1_1__leaf_net759),
    .X(net180));
 sky130_fd_sc_hd__mux4_1 c255 (.A0(net160),
    .A1(net60),
    .A2(net860),
    .A3(net943),
    .S0(net960),
    .S1(clknet_1_0__leaf_net901),
    .X(net910));
 sky130_fd_sc_hd__mux4_1 c256 (.A0(net47),
    .A1(clknet_1_0__leaf_net177),
    .A2(clknet_1_1__leaf_net924),
    .A3(clknet_1_0__leaf_net180),
    .S0(clknet_1_1__leaf_net910),
    .S1(clknet_1_0__leaf_net901),
    .X(net181));
 sky130_fd_sc_hd__mux4_1 c257 (.A0(net35),
    .A1(net62),
    .A2(net1038),
    .A3(net60),
    .S0(net1024),
    .S1(clknet_1_1__leaf_net901),
    .X(net182));
 sky130_fd_sc_hd__mux4_1 c258 (.A0(net59),
    .A1(clknet_1_0__leaf_net180),
    .A2(net884),
    .A3(net952),
    .S0(net52),
    .S1(clknet_1_1__leaf_net901),
    .X(net183));
 sky130_fd_sc_hd__mux4_1 c259 (.A0(clknet_1_1__leaf_net177),
    .A1(net1044),
    .A2(net29),
    .A3(net702),
    .S0(net899),
    .S1(clknet_1_1__leaf_net759),
    .X(net184));
 sky130_fd_sc_hd__mux4_2 c260 (.A0(net171),
    .A1(net58),
    .A2(net65),
    .A3(net173),
    .S0(net749),
    .S1(clknet_1_0__leaf_net759),
    .X(net185));
 sky130_fd_sc_hd__mux4_2 c261 (.A0(net1018),
    .A1(net185),
    .A2(net952),
    .A3(net749),
    .S0(clknet_1_0__leaf_net759),
    .S1(clknet_1_0__leaf_net901),
    .X(net186));
 sky130_fd_sc_hd__mux4_2 c262 (.A0(clknet_1_0__leaf_net186),
    .A1(net112),
    .A2(net854),
    .A3(net174),
    .S0(net749),
    .S1(clknet_1_0__leaf_net901),
    .X(net187));
 sky130_fd_sc_hd__mux4_2 c263 (.A0(clknet_1_0__leaf_net177),
    .A1(net187),
    .A2(clknet_1_1__leaf_net186),
    .A3(clknet_1_0__leaf_net905),
    .S0(net885),
    .S1(clknet_1_0__leaf_net759),
    .X(net188));
 sky130_fd_sc_hd__a21bo_1 c264 (.A1(net1024),
    .A2(net993),
    .B1_N(net980),
    .X(net189));
 sky130_fd_sc_hd__a21bo_2 c265 (.A1(net1016),
    .A2(net1003),
    .B1_N(net979),
    .X(net190));
 sky130_fd_sc_hd__a21bo_4 c266 (.A1(net998),
    .A2(net976),
    .B1_N(net1016),
    .X(net191));
 sky130_fd_sc_hd__a21bo_4 c267 (.A1(net977),
    .A2(net74),
    .B1_N(net998),
    .X(net192));
 sky130_fd_sc_hd__a41o_2 c268 (.A1(net81),
    .A2(net74),
    .A3(net191),
    .A4(net1009),
    .B1(net976),
    .X(net193));
 sky130_fd_sc_hd__a21bo_2 c269 (.A1(net980),
    .A2(net87),
    .B1_N(net976),
    .X(net194));
 sky130_fd_sc_hd__a41o_2 c270 (.A1(net1025),
    .A2(net75),
    .A3(net703),
    .A4(net977),
    .B1(net1005),
    .X(net195));
 sky130_fd_sc_hd__a21bo_2 c271 (.A1(net193),
    .A2(net703),
    .B1_N(net976),
    .X(net196));
 sky130_fd_sc_hd__a21bo_4 c272 (.A1(net827),
    .A2(net974),
    .B1_N(net976),
    .X(net197));
 sky130_fd_sc_hd__a21bo_2 c273 (.A1(net67),
    .A2(net191),
    .B1_N(net976),
    .X(net198));
 sky130_fd_sc_hd__a21bo_2 c274 (.A1(net193),
    .A2(net192),
    .B1_N(net984),
    .X(net199));
 sky130_fd_sc_hd__a41o_2 c275 (.A1(net974),
    .A2(net78),
    .A3(net191),
    .A4(net967),
    .B1(net976),
    .X(net200));
 sky130_fd_sc_hd__a31o_1 c276 (.A1(net196),
    .A2(net961),
    .A3(net68),
    .B1(net977),
    .X(net201));
 sky130_fd_sc_hd__a21bo_1 c277 (.A1(net1025),
    .A2(net974),
    .B1_N(net1014),
    .X(net202));
 sky130_fd_sc_hd__a21bo_1 c278 (.A1(net202),
    .A2(net198),
    .B1_N(net197),
    .X(net203));
 sky130_fd_sc_hd__a21bo_2 c279 (.A1(net201),
    .A2(net78),
    .B1_N(net963),
    .X(net204));
 sky130_fd_sc_hd__mux4_2 c280 (.A0(net192),
    .A1(net995),
    .A2(net974),
    .A3(net977),
    .S0(net196),
    .S1(net197),
    .X(net205));
 sky130_fd_sc_hd__mux4_2 c281 (.A0(net204),
    .A1(net202),
    .A2(net78),
    .A3(net967),
    .S0(net974),
    .S1(net963),
    .X(net206));
 sky130_fd_sc_hd__mux4_2 c282 (.A0(net1004),
    .A1(net197),
    .A2(net202),
    .A3(net963),
    .S0(net998),
    .S1(net976),
    .X(net207));
 sky130_fd_sc_hd__mux4_2 c283 (.A0(net194),
    .A1(net201),
    .A2(net703),
    .A3(net198),
    .S0(net963),
    .S1(net976),
    .X(net208));
 sky130_fd_sc_hd__mux4_2 c284 (.A0(net974),
    .A1(net205),
    .A2(net198),
    .A3(net204),
    .S0(net963),
    .S1(net976),
    .X(net209));
 sky130_fd_sc_hd__mux4_2 c285 (.A0(net208),
    .A1(net205),
    .A2(net209),
    .A3(net192),
    .S0(net974),
    .S1(net1004),
    .X(net210));
 sky130_fd_sc_hd__a21bo_2 c286 (.A1(net107),
    .A2(net840),
    .B1_N(net207),
    .X(net906));
 sky130_fd_sc_hd__a31o_4 c287 (.A1(net1023),
    .A2(net198),
    .A3(net1004),
    .B1(net853),
    .X(net211));
 sky130_fd_sc_hd__a31o_2 c288 (.A1(net1010),
    .A2(net208),
    .A3(net949),
    .B1(net206),
    .X(net917));
 sky130_fd_sc_hd__a31o_2 c289 (.A1(net194),
    .A2(net103),
    .A3(net962),
    .B1(net965),
    .X(net212));
 sky130_fd_sc_hd__a41o_4 c290 (.A1(net92),
    .A2(net87),
    .A3(net91),
    .A4(net1010),
    .B1(net977),
    .X(net213));
 sky130_fd_sc_hd__a41o_2 c291 (.A1(net90),
    .A2(net827),
    .A3(net967),
    .A4(net961),
    .B1(net106),
    .X(net214));
 sky130_fd_sc_hd__a21bo_1 c292 (.A1(net106),
    .A2(net944),
    .B1_N(net943),
    .X(net215));
 sky130_fd_sc_hd__a31o_1 c293 (.A1(net215),
    .A2(net214),
    .A3(net995),
    .B1(net933),
    .X(net216));
 sky130_fd_sc_hd__a21bo_4 c294 (.A1(net962),
    .A2(net104),
    .B1_N(net974),
    .X(net217));
 sky130_fd_sc_hd__a41o_2 c295 (.A1(net83),
    .A2(net1010),
    .A3(net991),
    .A4(net963),
    .B1(net213),
    .X(net218));
 sky130_fd_sc_hd__a31o_4 c296 (.A1(net944),
    .A2(net214),
    .A3(net213),
    .B1(net217),
    .X(net219));
 sky130_fd_sc_hd__a31o_2 c297 (.A1(net78),
    .A2(net853),
    .A3(net962),
    .B1(net208),
    .X(net220));
 sky130_fd_sc_hd__a41o_1 c298 (.A1(net213),
    .A2(net71),
    .A3(net96),
    .A4(net216),
    .B1(net944),
    .X(net221));
 sky130_fd_sc_hd__a31o_4 c299 (.A1(net832),
    .A2(net217),
    .A3(net219),
    .B1(net1025),
    .X(net222));
 sky130_fd_sc_hd__a31o_1 c300 (.A1(net222),
    .A2(net214),
    .A3(net936),
    .B1(net948),
    .X(net223));
 sky130_fd_sc_hd__a21bo_1 c301 (.A1(net222),
    .A2(net102),
    .B1_N(net950),
    .X(net224));
 sky130_fd_sc_hd__a31o_1 c302 (.A1(net86),
    .A2(net218),
    .A3(net219),
    .B1(net950),
    .X(net225));
 sky130_fd_sc_hd__a41o_1 c303 (.A1(net219),
    .A2(net224),
    .A3(net834),
    .A4(net950),
    .B1(net192),
    .X(net226));
 sky130_fd_sc_hd__mux4_2 c304 (.A0(net225),
    .A1(net213),
    .A2(net222),
    .A3(net1013),
    .S0(net96),
    .S1(net102),
    .X(net227));
 sky130_fd_sc_hd__mux4_1 c305 (.A0(net227),
    .A1(net832),
    .A2(net222),
    .A3(net950),
    .S0(net202),
    .S1(net962),
    .X(net228));
 sky130_fd_sc_hd__mux4_1 c306 (.A0(net102),
    .A1(net223),
    .A2(net933),
    .A3(net213),
    .S0(net962),
    .S1(net227),
    .X(net229));
 sky130_fd_sc_hd__mux4_1 c307 (.A0(net86),
    .A1(net227),
    .A2(net933),
    .A3(net202),
    .S0(net676),
    .S1(net988),
    .X(net230));
 sky130_fd_sc_hd__mux4_2 c308 (.A0(net71),
    .A1(net108),
    .A2(net193),
    .A3(net106),
    .S0(net984),
    .S1(net219),
    .X(net231));
 sky130_fd_sc_hd__a31o_1 c309 (.A1(net840),
    .A2(net104),
    .A3(net849),
    .B1(net1007),
    .X(net892));
 sky130_fd_sc_hd__a41o_4 c310 (.A1(net865),
    .A2(net123),
    .A3(net936),
    .A4(net1013),
    .B1(net1000),
    .X(net889));
 sky130_fd_sc_hd__mux4_1 c311 (.A0(net78),
    .A1(net120),
    .A2(net917),
    .A3(net119),
    .S0(net106),
    .S1(net941),
    .X(net232));
 sky130_fd_sc_hd__a31o_1 c312 (.A1(net191),
    .A2(net889),
    .A3(net1015),
    .B1(net941),
    .X(net233));
 sky130_fd_sc_hd__a31o_1 c313 (.A1(net233),
    .A2(net889),
    .A3(net960),
    .B1(net194),
    .X(net234));
 sky130_fd_sc_hd__a31o_1 c314 (.A1(net119),
    .A2(net79),
    .A3(net223),
    .X(net235));
 sky130_fd_sc_hd__a31o_4 c315 (.A1(net967),
    .A2(net118),
    .A3(net110),
    .B1(net127),
    .X(net236));
 sky130_fd_sc_hd__a41o_1 c316 (.A1(net108),
    .A2(net233),
    .A3(net218),
    .A4(net941),
    .B1(net745),
    .X(net237));
 sky130_fd_sc_hd__sdfbbn_2 c317 (.CLK_N(clknet_4_2_0_clk),
    .D(net118),
    .RESET_B(net227),
    .SCD(net125),
    .SCE(net889),
    .SET_B(net941),
    .Q(net239),
    .Q_N(net238));
 sky130_fd_sc_hd__a41o_1 c318 (.A1(net236),
    .A2(net73),
    .A3(net197),
    .A4(net1008),
    .B1(net745),
    .X(net240));
 sky130_fd_sc_hd__a41o_1 c319 (.A1(net225),
    .A2(net832),
    .A3(net996),
    .A4(net238),
    .B1(net745),
    .X(net241));
 sky130_fd_sc_hd__a41o_2 c320 (.A1(net91),
    .A2(net71),
    .A3(net840),
    .A4(net193),
    .B1(net110),
    .X(net242));
 sky130_fd_sc_hd__mux4_1 c321 (.A0(net127),
    .A1(net873),
    .A2(net233),
    .A3(net863),
    .S0(net242),
    .S1(net745),
    .X(net243));
 sky130_fd_sc_hd__a31o_1 c322 (.A1(net232),
    .A2(net233),
    .A3(net236),
    .B1(net209),
    .X(net244));
 sky130_fd_sc_hd__a41o_1 c323 (.A1(net221),
    .A2(net982),
    .A3(net126),
    .A4(net222),
    .B1(net727),
    .X(net245));
 sky130_fd_sc_hd__a31o_2 c324 (.A1(net847),
    .A2(net966),
    .A3(net684),
    .B1(net745),
    .X(net246));
 sky130_fd_sc_hd__mux4_2 c325 (.A0(net827),
    .A1(net239),
    .A2(net933),
    .A3(net246),
    .S0(net236),
    .S1(net727),
    .X(net247));
 sky130_fd_sc_hd__a41o_4 c326 (.A1(net247),
    .A2(net231),
    .A3(net849),
    .A4(net1),
    .B1(net699),
    .X(net248));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(net120),
    .A1(net248),
    .A2(net214),
    .A3(net238),
    .S0(net889),
    .S1(net236),
    .X(net249));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(net248),
    .A1(net238),
    .A2(net127),
    .A3(net242),
    .S0(net233),
    .S1(net721),
    .X(net250));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net121),
    .A1(net232),
    .A2(net248),
    .A3(net988),
    .S1(net727),
    .X(net251));
 sky130_fd_sc_hd__a41o_1 c330 (.A1(net1),
    .A2(net194),
    .A3(net248),
    .A4(net935),
    .B1(net79),
    .X(net252));
 sky130_fd_sc_hd__mux4_1 c331 (.A0(net109),
    .A1(net106),
    .A2(net248),
    .A3(net962),
    .S0(net868),
    .S1(net834),
    .X(net253));
 sky130_fd_sc_hd__a41o_1 c332 (.A1(net79),
    .A2(net1039),
    .A3(net1045),
    .A4(net842),
    .B1(net974),
    .X(net254));
 sky130_fd_sc_hd__mux4_1 c333 (.A0(net240),
    .A1(net142),
    .A2(net16),
    .A3(net101),
    .S0(net827),
    .S1(net761),
    .X(net255));
 sky130_fd_sc_hd__a41o_1 c334 (.A1(net223),
    .A2(net129),
    .A3(net240),
    .A4(net935),
    .B1(net760),
    .X(net256));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(net1039),
    .A1(net917),
    .A2(net198),
    .A3(net82),
    .S0(net1023),
    .S1(net664),
    .X(net257));
 sky130_fd_sc_hd__mux4_1 c336 (.A0(net214),
    .A1(net1039),
    .A2(net941),
    .A3(net677),
    .S0(net721),
    .S1(net761),
    .X(net258));
 sky130_fd_sc_hd__mux4_1 c337 (.A0(net104),
    .A1(net991),
    .A2(net198),
    .A3(net857),
    .S0(net721),
    .S1(net761),
    .X(net259));
 sky130_fd_sc_hd__mux4_1 c338 (.A0(net254),
    .A1(net1010),
    .A2(net1),
    .A3(net935),
    .S0(net79),
    .S1(net145),
    .X(net260));
 sky130_fd_sc_hd__mux4_2 c339 (.A0(net257),
    .A1(net19),
    .A2(net1012),
    .A3(net823),
    .S0(net664),
    .S1(net989),
    .X(net261));
 sky130_fd_sc_hd__mux4_2 c340 (.A0(net214),
    .A1(net212),
    .A2(net962),
    .A3(net257),
    .S0(net19),
    .S1(net714),
    .X(net262));
 sky130_fd_sc_hd__a41o_2 c341 (.A1(net1002),
    .A2(net1026),
    .A3(net867),
    .A4(net10),
    .B1(net899),
    .X(net263));
 sky130_fd_sc_hd__mux4_2 c342 (.A0(net86),
    .A1(net254),
    .A2(net891),
    .A3(net257),
    .S0(net958),
    .S1(net760),
    .X(net264));
 sky130_fd_sc_hd__mux4_1 c343 (.A0(net132),
    .A1(net967),
    .A2(net264),
    .A3(net130),
    .S0(net664),
    .S1(net677),
    .X(net265));
 sky130_fd_sc_hd__mux4_2 c344 (.A0(net123),
    .A1(net262),
    .A2(net1018),
    .A3(net261),
    .S0(net989),
    .S1(net732),
    .X(net266));
 sky130_fd_sc_hd__a41o_2 c345 (.A1(net123),
    .A2(net891),
    .A3(net259),
    .A4(net139),
    .B1(net721),
    .X(net267));
 sky130_fd_sc_hd__mux4_2 c346 (.A0(net123),
    .A1(net259),
    .A2(net207),
    .A3(net677),
    .S0(net745),
    .S1(net760),
    .X(net268));
 sky130_fd_sc_hd__mux4_2 c347 (.A0(net198),
    .A1(net109),
    .A2(net267),
    .A3(net941),
    .S0(net264),
    .S1(net899),
    .X(net269));
 sky130_fd_sc_hd__mux4_2 c348 (.A0(net259),
    .A1(net109),
    .A2(net254),
    .A3(net121),
    .S0(net857),
    .S1(net899),
    .X(net270));
 sky130_fd_sc_hd__mux4_2 c349 (.A0(net130),
    .A1(net1013),
    .A2(net270),
    .A3(net267),
    .S0(net258),
    .S1(net714),
    .X(net271));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(net258),
    .A1(net240),
    .A2(net262),
    .A3(net86),
    .S0(net958),
    .S1(net271),
    .X(net272));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net264),
    .A1(net270),
    .A2(net936),
    .A3(net132),
    .S0(net664),
    .S1(net1059),
    .X(net273));
 sky130_fd_sc_hd__mux4_1 c352 (.A0(net135),
    .A1(net248),
    .A2(net271),
    .A3(net973),
    .S0(net961),
    .S1(net760),
    .X(net274));
 sky130_fd_sc_hd__mux4_1 c353 (.A0(net39),
    .A1(net823),
    .A2(net42),
    .A3(net129),
    .S0(net212),
    .S1(net731),
    .X(net275));
 sky130_fd_sc_hd__mux4_1 c354 (.A0(clknet_1_0__leaf_net170),
    .A1(net857),
    .A2(net992),
    .A3(net823),
    .S0(net957),
    .S1(clknet_1_0__leaf_net758),
    .X(net276));
 sky130_fd_sc_hd__mux4_1 c355 (.A0(net40),
    .A1(net831),
    .A2(net865),
    .A3(net269),
    .S0(net264),
    .S1(net942),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 c356 (.A0(net152),
    .A1(net246),
    .A2(net264),
    .A3(net972),
    .S0(clknet_1_1__leaf_net170),
    .S1(net734),
    .X(net916));
 sky130_fd_sc_hd__mux4_1 c357 (.A0(net246),
    .A1(net152),
    .A2(net82),
    .A3(net865),
    .S0(net731),
    .S1(net762),
    .X(net278));
 sky130_fd_sc_hd__mux4_1 c358 (.A0(net42),
    .A1(net134),
    .A2(net868),
    .A3(net856),
    .S0(net1006),
    .S1(net1069),
    .X(net279));
 sky130_fd_sc_hd__mux4_2 c359 (.A0(net1040),
    .A1(net134),
    .A2(net993),
    .A3(net1024),
    .S0(net955),
    .S1(net1008),
    .X(net923));
 sky130_fd_sc_hd__mux4_1 c360 (.A0(net966),
    .A1(net962),
    .A2(net866),
    .A3(net891),
    .S0(net955),
    .S1(net944),
    .X(net280));
 sky130_fd_sc_hd__mux4_1 c361 (.A0(net33),
    .A1(net280),
    .A2(net1004),
    .A3(net955),
    .S0(clknet_1_0__leaf_net758),
    .S1(net762),
    .X(net281));
 sky130_fd_sc_hd__mux4_1 c362 (.A0(net858),
    .A1(net275),
    .A2(net193),
    .A3(net279),
    .S0(net955),
    .S1(net1048),
    .X(net282));
 sky130_fd_sc_hd__mux4_1 c363 (.A0(net37),
    .A1(net152),
    .A2(net1011),
    .A3(net955),
    .S0(net271),
    .S1(net930),
    .X(net283));
 sky130_fd_sc_hd__mux4_2 c364 (.A0(net150),
    .A1(net225),
    .A2(net993),
    .A3(net1000),
    .S0(net955),
    .S1(net872),
    .X(net284));
 sky130_fd_sc_hd__mux4_1 c365 (.A0(net193),
    .A1(net1012),
    .A2(net955),
    .A3(net713),
    .S0(clknet_1_0__leaf_net758),
    .S1(net920),
    .X(net285));
 sky130_fd_sc_hd__mux4_1 c366 (.A0(clknet_1_0__leaf_net276),
    .A1(net39),
    .A2(net889),
    .A3(net1011),
    .S0(net943),
    .S1(net721),
    .X(net286));
 sky130_fd_sc_hd__mux4_1 c367 (.A0(net1031),
    .A1(net150),
    .A2(net844),
    .A3(net1040),
    .S0(net692),
    .S1(net713),
    .X(net287));
 sky130_fd_sc_hd__mux4_1 c368 (.A0(net142),
    .A1(net285),
    .A2(net955),
    .A3(net944),
    .S0(net756),
    .S1(net763),
    .X(net288));
 sky130_fd_sc_hd__a41o_1 c369 (.A1(net121),
    .A2(net955),
    .A3(net275),
    .A4(net692),
    .B1(net764),
    .X(net918));
 sky130_fd_sc_hd__mux4_1 c370 (.A0(net205),
    .A1(net837),
    .A2(net918),
    .A3(net955),
    .S0(net925),
    .S1(net764),
    .X(net912));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(clknet_1_1__leaf_net281),
    .A1(net918),
    .A2(net40),
    .A3(net30),
    .S0(net731),
    .S1(net764),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net1032),
    .A1(net31),
    .A2(net923),
    .A3(net247),
    .S0(net713),
    .S1(net1056),
    .X(net290));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net289),
    .A1(net263),
    .A2(net956),
    .A3(net39),
    .S0(net1006),
    .S1(net764),
    .X(net911));
 sky130_fd_sc_hd__mux4_1 c374 (.A0(net145),
    .A1(clknet_1_1__leaf_net902),
    .A2(net271),
    .A3(net834),
    .S0(net134),
    .S1(net702),
    .X(net291));
 sky130_fd_sc_hd__mux4_1 c375 (.A0(net66),
    .A1(net856),
    .A2(net1006),
    .A3(clknet_1_0__leaf_net179),
    .S0(net974),
    .S1(net952),
    .X(net292));
 sky130_fd_sc_hd__mux4_1 c376 (.A0(net49),
    .A1(net134),
    .A2(net1079),
    .A3(net888),
    .S0(net997),
    .S1(net1015),
    .X(net293));
 sky130_fd_sc_hd__mux4_1 c377 (.A0(net50),
    .A1(net880),
    .A2(net162),
    .A3(clknet_1_1__leaf_net177),
    .S0(net1013),
    .S1(net702),
    .X(net294));
 sky130_fd_sc_hd__mux4_1 c378 (.A0(net271),
    .A1(clknet_1_1__leaf_net180),
    .A2(net960),
    .A3(net898),
    .S0(net997),
    .S1(net925),
    .X(net295));
 sky130_fd_sc_hd__mux4_1 c379 (.A0(net262),
    .A1(net56),
    .A2(net975),
    .A3(net992),
    .S0(net752),
    .S1(clknet_1_1__leaf_net901),
    .X(net296));
 sky130_fd_sc_hd__mux4_1 c380 (.A0(net264),
    .A1(net981),
    .A2(net992),
    .A3(net844),
    .S0(net972),
    .S1(net927),
    .X(net297));
 sky130_fd_sc_hd__mux4_1 c381 (.A0(net868),
    .A1(net297),
    .A2(net271),
    .A3(net952),
    .S0(net899),
    .S1(net748),
    .X(net298));
 sky130_fd_sc_hd__mux4_1 c382 (.A0(net53),
    .A1(net31),
    .A2(net889),
    .A3(net65),
    .S0(clknet_1_1__leaf_net759),
    .S1(net765),
    .X(net299));
 sky130_fd_sc_hd__mux4_1 c383 (.A0(net1024),
    .A1(net270),
    .A2(net1037),
    .A3(net1007),
    .S0(net65),
    .S1(net992),
    .X(net300));
 sky130_fd_sc_hd__mux4_1 c384 (.A0(net300),
    .A1(net913),
    .A2(net1038),
    .A3(net284),
    .S0(clknet_1_1__leaf_net709),
    .S1(net748),
    .X(net301));
 sky130_fd_sc_hd__mux4_1 c385 (.A0(clknet_1_1__leaf_net179),
    .A1(net972),
    .A2(net904),
    .A3(net954),
    .S0(net752),
    .S1(net766),
    .X(net302));
 sky130_fd_sc_hd__mux4_1 c386 (.A0(net302),
    .A1(net31),
    .A2(net1021),
    .A3(net880),
    .S0(net697),
    .S1(net763),
    .X(net303));
 sky130_fd_sc_hd__mux4_1 c387 (.A0(net1079),
    .A1(net264),
    .A2(net952),
    .A3(net975),
    .S0(net897),
    .S1(net765),
    .X(net304));
 sky130_fd_sc_hd__mux4_1 c388 (.A0(net299),
    .A1(net952),
    .A2(net37),
    .A3(net997),
    .S0(net749),
    .S1(net766),
    .X(net305));
 sky130_fd_sc_hd__mux4_1 c389 (.A0(net975),
    .A1(net825),
    .A2(net139),
    .A3(net748),
    .S0(net752),
    .S1(clknet_1_1__leaf_net759),
    .X(net306));
 sky130_fd_sc_hd__mux4_1 c390 (.A0(net52),
    .A1(net972),
    .A2(net952),
    .A3(net702),
    .S0(net762),
    .S1(net765),
    .X(net307));
 sky130_fd_sc_hd__mux4_1 c391 (.A0(net307),
    .A1(net66),
    .A2(net888),
    .A3(net990),
    .S0(net897),
    .S1(net766),
    .X(net308));
 sky130_fd_sc_hd__mux4_2 c392 (.A0(net58),
    .A1(net52),
    .A2(net825),
    .A3(net954),
    .S0(net271),
    .S1(net766),
    .X(net309));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net308),
    .A1(net306),
    .A2(net66),
    .A3(net975),
    .S0(net952),
    .S1(net1023),
    .X(net310));
 sky130_fd_sc_hd__mux4_1 c394 (.A0(net293),
    .A1(net1021),
    .A2(net856),
    .A3(net919),
    .S0(net975),
    .S1(clknet_1_1__leaf_net744),
    .X(net311));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net292),
    .A1(net310),
    .A2(net37),
    .A3(net975),
    .S0(net748),
    .S1(net765),
    .X(net312));
 sky130_fd_sc_hd__xnor2_4 c396 (.A(net1012),
    .B(net204),
    .Y(net313));
 sky130_fd_sc_hd__a21bo_2 c397 (.A1(net81),
    .A2(net205),
    .B1_N(net963),
    .X(net314));
 sky130_fd_sc_hd__a41o_2 c398 (.A1(net984),
    .A2(net85),
    .A3(net314),
    .A4(net191),
    .B1(net963),
    .X(net315));
 sky130_fd_sc_hd__xnor2_2 c399 (.A(net313),
    .B(net1005),
    .Y(net316));
 sky130_fd_sc_hd__a21bo_2 c400 (.A1(net996),
    .A2(net75),
    .B1_N(net192),
    .X(net317));
 sky130_fd_sc_hd__a21bo_2 c401 (.A1(net703),
    .A2(net316),
    .B1_N(net964),
    .X(net318));
 sky130_fd_sc_hd__a21bo_1 c402 (.A1(net318),
    .A2(net968),
    .B1_N(net967),
    .X(net319));
 sky130_fd_sc_hd__a21bo_1 c403 (.A1(net1009),
    .A2(net1022),
    .B1_N(net313),
    .X(net900));
 sky130_fd_sc_hd__a41o_2 c404 (.A1(net1021),
    .A2(net996),
    .A3(net74),
    .A4(net968),
    .B1(net945),
    .X(net320));
 sky130_fd_sc_hd__a21bo_4 c405 (.A1(net968),
    .A2(net318),
    .B1_N(net945),
    .X(net321));
 sky130_fd_sc_hd__a41o_2 c406 (.A1(net320),
    .A2(net314),
    .A3(net945),
    .A4(net967),
    .B1(net996),
    .X(net322));
 sky130_fd_sc_hd__a41o_2 c407 (.A1(net1005),
    .A2(net939),
    .A3(net963),
    .A4(net945),
    .B1(net1022),
    .X(net323));
 sky130_fd_sc_hd__a21bo_4 c408 (.A1(net961),
    .A2(net321),
    .B1_N(net945),
    .X(net324));
 sky130_fd_sc_hd__mux4_2 c409 (.A0(net315),
    .A1(net209),
    .A2(net321),
    .A3(net322),
    .S0(net1009),
    .S1(net945),
    .X(net325));
 sky130_fd_sc_hd__mux4_2 c410 (.A0(net74),
    .A1(net322),
    .A2(net321),
    .A3(net968),
    .S0(net324),
    .S1(net945),
    .X(net326));
 sky130_fd_sc_hd__mux4_2 c411 (.A0(net939),
    .A1(net326),
    .A2(net318),
    .A3(net324),
    .S0(net321),
    .S1(net1012),
    .X(net327));
 sky130_fd_sc_hd__mux4_2 c412 (.A0(net323),
    .A1(net325),
    .A2(net320),
    .A3(net207),
    .S0(net967),
    .S1(net945),
    .X(net328));
 sky130_fd_sc_hd__a21bo_4 c413 (.A1(net327),
    .A2(net1006),
    .B1_N(net946),
    .X(net929));
 sky130_fd_sc_hd__mux4_2 c414 (.A0(net321),
    .A1(net929),
    .A2(net314),
    .A3(net328),
    .S0(net196),
    .S1(net967),
    .X(net329));
 sky130_fd_sc_hd__mux4_2 c415 (.A0(net201),
    .A1(net328),
    .A2(net329),
    .A3(net322),
    .S0(net318),
    .S1(net945),
    .X(net330));
 sky130_fd_sc_hd__a41o_1 c416 (.A1(net329),
    .A2(net206),
    .A3(net946),
    .A4(net996),
    .B1(net328),
    .X(net331));
 sky130_fd_sc_hd__mux4_1 c417 (.A0(net204),
    .A1(net326),
    .A2(net206),
    .A3(net331),
    .S0(net322),
    .S1(net945),
    .X(net332));
 sky130_fd_sc_hd__a41o_1 c418 (.A1(net75),
    .A2(net836),
    .A3(net313),
    .A4(net1025),
    .B1(net327),
    .X(net333));
 sky130_fd_sc_hd__dlymetal6s2s_1 c419 (.A(net663),
    .X(net334));
 sky130_fd_sc_hd__a21bo_1 c420 (.A1(net949),
    .A2(net207),
    .B1_N(net965),
    .X(net335));
 sky130_fd_sc_hd__a21bo_2 c421 (.A1(net91),
    .A2(net313),
    .B1_N(net984),
    .X(net926));
 sky130_fd_sc_hd__a21bo_1 c422 (.A1(net320),
    .A2(net996),
    .B1_N(net222),
    .X(net336));
 sky130_fd_sc_hd__a41o_1 c423 (.A1(net334),
    .A2(net1025),
    .A3(net213),
    .A4(net1022),
    .B1(net75),
    .X(net337));
 sky130_fd_sc_hd__a31o_4 c424 (.A1(net836),
    .A2(net320),
    .A3(net926),
    .B1(net998),
    .X(net338));
 sky130_fd_sc_hd__a21bo_1 c425 (.A1(net200),
    .A2(net333),
    .B1_N(net99),
    .X(net339));
 sky130_fd_sc_hd__mux4_1 c426 (.A0(net80),
    .A1(net337),
    .A2(net192),
    .A3(net335),
    .S0(net320),
    .S1(net963),
    .X(net340));
 sky130_fd_sc_hd__buf_1 c427 (.A(net663),
    .X(net341));
 sky130_fd_sc_hd__a41o_2 c428 (.A1(net216),
    .A2(net93),
    .A3(net313),
    .A4(net962),
    .B1(net965),
    .X(net342));
 sky130_fd_sc_hd__a41o_2 c429 (.A1(net202),
    .A2(net327),
    .A3(net337),
    .A4(net192),
    .B1(net99),
    .X(net343));
 sky130_fd_sc_hd__a31o_1 c430 (.A1(net103),
    .A2(net937),
    .A3(net224),
    .B1(net341),
    .X(net344));
 sky130_fd_sc_hd__a41o_2 c431 (.A1(net1021),
    .A2(net937),
    .A3(net103),
    .A4(net338),
    .B1(net341),
    .X(net345));
 sky130_fd_sc_hd__sdfbbn_2 c432 (.CLK_N(clknet_4_8_0_clk),
    .D(net325),
    .RESET_B(net342),
    .SCD(net948),
    .SCE(net338),
    .SET_B(net321),
    .Q(net347),
    .Q_N(net346));
 sky130_fd_sc_hd__a21bo_1 c433 (.A1(net337),
    .A2(net347),
    .B1_N(net846),
    .X(net348));
 sky130_fd_sc_hd__a41o_1 c434 (.A1(net335),
    .A2(net221),
    .A3(net948),
    .A4(net1052),
    .B1(net937),
    .X(net349));
 sky130_fd_sc_hd__a41o_2 c435 (.A1(net339),
    .A2(net937),
    .A3(net968),
    .A4(net663),
    .B1(net698),
    .X(net350));
 sky130_fd_sc_hd__a41o_1 c436 (.A1(net853),
    .A2(net348),
    .A3(net336),
    .A4(net937),
    .B1(net1061),
    .X(net351));
 sky130_fd_sc_hd__a41o_1 c437 (.A1(net341),
    .A2(net980),
    .A3(net937),
    .A4(net939),
    .B1(net663),
    .X(net352));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(net338),
    .A1(net348),
    .A2(net946),
    .A3(net346),
    .S0(net937),
    .S1(net337),
    .X(net353));
 sky130_fd_sc_hd__mux4_2 c439 (.A0(net353),
    .A1(net348),
    .A2(net213),
    .A3(net937),
    .S0(net209),
    .S1(net1009),
    .X(net354));
 sky130_fd_sc_hd__mux4_1 c440 (.A0(net231),
    .A1(net127),
    .A2(net993),
    .A3(net947),
    .S0(net941),
    .S1(net988),
    .X(net355));
 sky130_fd_sc_hd__mux4_1 c441 (.A0(net355),
    .A1(net125),
    .A2(net1005),
    .A3(net998),
    .S0(net842),
    .S1(net1054),
    .X(net356));
 sky130_fd_sc_hd__mux4_1 c442 (.A0(net197),
    .A1(net126),
    .A2(net247),
    .A3(net354),
    .S0(net74),
    .S1(net937),
    .X(net357));
 sky130_fd_sc_hd__mux4_1 c443 (.A0(net127),
    .A1(net219),
    .A2(net325),
    .A3(net236),
    .S0(net209),
    .S1(net231),
    .X(net358));
 sky130_fd_sc_hd__mux4_2 c444 (.A0(net994),
    .A1(net338),
    .A2(net103),
    .A3(net339),
    .S0(net978),
    .S1(net655),
    .X(net359));
 sky130_fd_sc_hd__mux4_2 c445 (.A0(net938),
    .A1(net982),
    .A2(net950),
    .A3(net961),
    .S0(net699),
    .S1(net727),
    .X(net360));
 sky130_fd_sc_hd__mux4_1 c446 (.A0(net99),
    .A1(net126),
    .A2(net227),
    .A3(net350),
    .S0(net345),
    .S1(net727),
    .X(net361));
 sky130_fd_sc_hd__mux4_2 c447 (.A0(net208),
    .A1(net321),
    .A2(net949),
    .A3(net190),
    .S0(net75),
    .S1(net217),
    .X(net890));
 sky130_fd_sc_hd__mux4_1 c448 (.A0(net950),
    .A1(net355),
    .A2(net350),
    .A3(net236),
    .S0(net983),
    .S1(net218),
    .X(net362));
 sky130_fd_sc_hd__mux4_1 c449 (.A0(net358),
    .A1(net343),
    .A2(net926),
    .A3(net350),
    .S0(net890),
    .S1(net222),
    .X(net363));
 sky130_fd_sc_hd__mux4_2 c450 (.A0(net75),
    .A1(net994),
    .A2(net91),
    .A3(net993),
    .S0(net346),
    .S1(net948),
    .X(net364));
 sky130_fd_sc_hd__mux4_1 c451 (.A0(net242),
    .A1(net338),
    .A2(net247),
    .A3(net354),
    .S0(net965),
    .S1(net937),
    .X(net365));
 sky130_fd_sc_hd__mux4_1 c452 (.A0(net939),
    .A1(net889),
    .A2(net365),
    .A3(net988),
    .S0(net730),
    .S1(net770),
    .X(net366));
 sky130_fd_sc_hd__sdfbbp_1 c453 (.CLK(clknet_4_9_0_clk),
    .D(net354),
    .RESET_B(net91),
    .SCD(net342),
    .SCE(net358),
    .SET_B(net730),
    .Q(net368),
    .Q_N(net367));
 sky130_fd_sc_hd__mux4_1 c454 (.A0(net365),
    .A1(net359),
    .A2(net1016),
    .A3(net1003),
    .S0(net730),
    .S1(net987),
    .X(net369));
 sky130_fd_sc_hd__mux4_1 c455 (.A0(net336),
    .A1(net325),
    .A2(net365),
    .A3(net676),
    .S0(net698),
    .S1(net1057),
    .X(net370));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(net364),
    .A1(net890),
    .A2(net1008),
    .A3(net222),
    .S0(net994),
    .S1(net1067),
    .X(net371));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(net873),
    .A1(net336),
    .A2(net1022),
    .A3(net371),
    .S0(net1054),
    .S1(net1050),
    .X(net372));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(net246),
    .A1(net0),
    .A2(net371),
    .A3(net994),
    .S0(net654),
    .S1(net1065),
    .X(net373));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net206),
    .A1(net350),
    .A2(net365),
    .A3(net359),
    .S0(net771),
    .S1(net773),
    .X(net374));
 sky130_fd_sc_hd__mux4_2 c460 (.A0(net197),
    .A1(net238),
    .A2(net933),
    .A3(net654),
    .S0(net699),
    .S1(net773),
    .X(net375));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net371),
    .A1(net222),
    .A2(net375),
    .A3(net242),
    .S0(net772),
    .S1(net773),
    .X(net376));
 sky130_fd_sc_hd__mux4_1 c462 (.A0(net996),
    .A1(net190),
    .A2(net1000),
    .A3(net926),
    .S0(net1042),
    .S1(net655),
    .X(net377));
 sky130_fd_sc_hd__mux4_1 c463 (.A0(net377),
    .A1(net938),
    .A2(net268),
    .A3(net891),
    .S0(net247),
    .S1(net774),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 c464 (.A0(net948),
    .A1(net984),
    .A2(net367),
    .A3(net735),
    .S0(net745),
    .S1(net771),
    .X(net379));
 sky130_fd_sc_hd__mux4_1 c465 (.A0(net368),
    .A1(net1043),
    .A2(net239),
    .A3(net940),
    .S0(net359),
    .S1(net966),
    .X(net380));
 sky130_fd_sc_hd__mux4_1 c466 (.A0(net227),
    .A1(net324),
    .A2(net125),
    .A3(net938),
    .S0(net1016),
    .S1(net774),
    .X(net381));
 sky130_fd_sc_hd__mux4_1 c467 (.A0(net131),
    .A1(net938),
    .A2(net979),
    .A3(net994),
    .S0(net989),
    .S1(net767),
    .X(net382));
 sky130_fd_sc_hd__mux4_1 c468 (.A0(net359),
    .A1(net350),
    .A2(net227),
    .A3(net953),
    .S0(net958),
    .S1(net988),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 c469 (.A0(net81),
    .A1(net872),
    .A2(net997),
    .A3(net1003),
    .S0(net994),
    .S1(net772),
    .X(net384));
 sky130_fd_sc_hd__mux4_1 c470 (.A0(net870),
    .A1(net378),
    .A2(net1042),
    .A3(net267),
    .S0(net0),
    .S1(net984),
    .X(net385));
 sky130_fd_sc_hd__mux4_1 c471 (.A0(net129),
    .A1(net239),
    .A2(net81),
    .A3(net323),
    .S0(net270),
    .S1(net217),
    .X(net386));
 sky130_fd_sc_hd__mux4_1 c472 (.A0(net936),
    .A1(net386),
    .A2(net890),
    .A3(net1000),
    .S0(net684),
    .S1(net988),
    .X(net387));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(net261),
    .A1(net387),
    .A2(net263),
    .A3(net948),
    .S0(net676),
    .S1(clknet_1_1__leaf_net775),
    .X(net388));
 sky130_fd_sc_hd__mux4_1 c474 (.A0(net360),
    .A1(net263),
    .A2(net684),
    .A3(net729),
    .S0(net767),
    .S1(clknet_1_0__leaf_net777),
    .X(net389));
 sky130_fd_sc_hd__mux4_1 c475 (.A0(net131),
    .A1(net948),
    .A2(net270),
    .A3(net1021),
    .S0(net988),
    .S1(clknet_1_0__leaf_net777),
    .X(net390));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(net190),
    .A1(net1008),
    .A2(net984),
    .A3(net382),
    .S0(net933),
    .S1(clknet_1_1__leaf_net777),
    .X(net391));
 sky130_fd_sc_hd__mux4_2 c477 (.A0(net938),
    .A1(net961),
    .A2(net841),
    .A3(net1008),
    .S0(net994),
    .S1(net940),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(net321),
    .A1(net327),
    .A2(clknet_1_0__leaf_net389),
    .A3(net343),
    .S0(net116),
    .S1(net103),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(net386),
    .A1(net387),
    .A2(net74),
    .A3(net392),
    .S0(net378),
    .S1(net729),
    .X(net394));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net393),
    .A1(net222),
    .A2(clknet_1_0__leaf_net389),
    .A3(net368),
    .S0(net732),
    .S1(net778),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net384),
    .A1(net382),
    .A2(net360),
    .A3(net948),
    .S0(net392),
    .S1(net779),
    .X(net396));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(net387),
    .A1(net938),
    .A2(net947),
    .A3(net396),
    .S0(net979),
    .S1(net779),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net23),
    .A1(net74),
    .A2(net392),
    .A3(clknet_1_0__leaf_net710),
    .S0(clknet_1_0__leaf_net777),
    .S1(net778),
    .X(net398));
 sky130_fd_sc_hd__mux4_1 c484 (.A0(net279),
    .A1(net837),
    .A2(net849),
    .A3(net1037),
    .S0(net1048),
    .S1(net1055),
    .X(net399));
 sky130_fd_sc_hd__mux4_1 c485 (.A0(net382),
    .A1(net360),
    .A2(net116),
    .A3(clknet_1_0__leaf_net398),
    .S0(net270),
    .S1(net767),
    .X(net400));
 sky130_fd_sc_hd__mux4_1 c486 (.A0(net343),
    .A1(net866),
    .A2(net269),
    .A3(net30),
    .S0(net246),
    .S1(net779),
    .X(net401));
 sky130_fd_sc_hd__mux4_1 c487 (.A0(net266),
    .A1(net919),
    .A2(clknet_1_0__leaf_net911),
    .A3(net956),
    .S0(net912),
    .S1(net246),
    .X(net402));
 sky130_fd_sc_hd__mux4_1 c488 (.A0(net333),
    .A1(net116),
    .A2(net343),
    .A3(net1019),
    .S0(net236),
    .S1(net729),
    .X(net403));
 sky130_fd_sc_hd__mux4_1 c489 (.A0(clknet_1_1__leaf_net276),
    .A1(clknet_1_1__leaf_net389),
    .A2(net863),
    .A3(net30),
    .S0(net691),
    .S1(net921),
    .X(net404));
 sky130_fd_sc_hd__mux4_1 c490 (.A0(net218),
    .A1(net10),
    .A2(net345),
    .A3(net266),
    .S0(net343),
    .S1(net987),
    .X(net405));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(net403),
    .A1(net926),
    .A2(net248),
    .A3(net247),
    .S0(net691),
    .S1(net757),
    .X(net406));
 sky130_fd_sc_hd__mux4_1 c492 (.A0(net390),
    .A1(net849),
    .A2(net1008),
    .A3(net923),
    .S0(net997),
    .S1(net782),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(net837),
    .A1(net919),
    .A2(net30),
    .A3(net1023),
    .S0(net1006),
    .S1(net675),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(net891),
    .A1(net931),
    .A2(clknet_1_1__leaf_net758),
    .A3(net771),
    .S0(net783),
    .S1(net784),
    .X(net409));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(clknet_1_0__leaf_net281),
    .A1(clknet_1_0__leaf_net276),
    .A2(net125),
    .A3(net983),
    .S0(net1038),
    .S1(net784),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(net284),
    .A1(net266),
    .A2(net942),
    .A3(net116),
    .S0(net724),
    .S1(net767),
    .X(net411));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net116),
    .A1(net1019),
    .A2(net248),
    .A3(net908),
    .S0(net989),
    .S1(net784),
    .X(net412));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(net890),
    .A1(net267),
    .A2(net139),
    .A3(net725),
    .S0(net783),
    .S1(net784),
    .X(net413));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(net30),
    .A1(net956),
    .A2(clknet_1_0__leaf_net398),
    .A3(net723),
    .S0(net757),
    .S1(net784),
    .X(net414));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(net360),
    .A1(net1006),
    .A2(net1027),
    .A3(net725),
    .S0(net780),
    .S1(net784),
    .X(net415));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(net395),
    .A1(net923),
    .A2(net415),
    .A3(net982),
    .S0(net30),
    .S1(net782),
    .X(net416));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(net953),
    .A1(net922),
    .A2(net16),
    .A3(net724),
    .S0(net780),
    .S1(net784),
    .X(net417));
 sky130_fd_sc_hd__mux4_2 c503 (.A0(net125),
    .A1(net417),
    .A2(net918),
    .A3(net15),
    .S0(net36),
    .S1(net782),
    .X(net418));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net414),
    .A1(net904),
    .A2(net942),
    .A3(net1019),
    .S0(net761),
    .S1(net767),
    .X(net419));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(net419),
    .A1(net982),
    .A2(net324),
    .A3(net129),
    .S0(net30),
    .S1(net757),
    .X(net420));
 sky130_fd_sc_hd__mux4_1 c526 (.A0(net350),
    .A1(net992),
    .A2(net894),
    .A3(net908),
    .S0(net920),
    .S1(net784),
    .X(net421));
 sky130_fd_sc_hd__mux4_1 c527 (.A0(net834),
    .A1(net284),
    .A2(net312),
    .A3(net304),
    .S0(net894),
    .S1(clknet_1_1__leaf_net901),
    .X(net422));
 sky130_fd_sc_hd__buf_1 c528 (.A(net690),
    .X(net423));
 sky130_fd_sc_hd__a31o_1 c529 (.A1(net87),
    .A2(net331),
    .A3(net1019),
    .B1(net999),
    .X(net424));
 sky130_fd_sc_hd__a21bo_1 c530 (.A1(net318),
    .A2(net197),
    .B1_N(net929),
    .X(net425));
 sky130_fd_sc_hd__a41o_2 c531 (.A1(net197),
    .A2(net324),
    .A3(net964),
    .A4(net999),
    .B1(net1022),
    .X(net426));
 sky130_fd_sc_hd__a41o_2 c532 (.A1(net328),
    .A2(net314),
    .A3(net969),
    .A4(net426),
    .B1(net980),
    .X(net427));
 sky130_fd_sc_hd__a31o_1 c533 (.A1(net323),
    .A2(net939),
    .A3(net68),
    .B1(net672),
    .X(net428));
 sky130_fd_sc_hd__a21bo_2 c534 (.A1(net427),
    .A2(net948),
    .B1_N(net980),
    .X(net429));
 sky130_fd_sc_hd__a21bo_1 c535 (.A1(net85),
    .A2(net209),
    .B1_N(net1014),
    .X(net430));
 sky130_fd_sc_hd__a31o_1 c536 (.A1(net425),
    .A2(net318),
    .A3(net939),
    .B1(net964),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_1 c537 (.A(net690),
    .X(net432));
 sky130_fd_sc_hd__a21bo_1 c538 (.A1(net1016),
    .A2(net318),
    .B1_N(net994),
    .X(net433));
 sky130_fd_sc_hd__mux4_2 c539 (.A0(net948),
    .A1(net200),
    .A2(net1009),
    .A3(net425),
    .S0(net192),
    .S1(net426),
    .X(net434));
 sky130_fd_sc_hd__sdfrbp_1 c540 (.CLK(clknet_4_8_0_clk),
    .D(net434),
    .RESET_B(net87),
    .SCD(net433),
    .SCE(net946),
    .Q(net436),
    .Q_N(net435));
 sky130_fd_sc_hd__a41o_4 c541 (.A1(net430),
    .A2(net1025),
    .A3(net426),
    .A4(net969),
    .B1(net429),
    .X(net437));
 sky130_fd_sc_hd__sdfbbn_2 c542 (.CLK_N(clknet_4_8_0_clk),
    .D(net433),
    .RESET_B(net969),
    .SCD(net423),
    .SCE(net85),
    .SET_B(net434),
    .Q(net915),
    .Q_N(net438));
 sky130_fd_sc_hd__sdfbbn_2 c543 (.CLK_N(clknet_4_10_0_clk),
    .D(net1062),
    .RESET_B(net314),
    .SCD(net435),
    .SCE(net87),
    .SET_B(net434),
    .Q(net907),
    .Q_N(net439));
 sky130_fd_sc_hd__a41o_1 c544 (.A1(net431),
    .A2(net437),
    .A3(net969),
    .A4(net1060),
    .B1(net439),
    .X(net440));
 sky130_fd_sc_hd__a41o_1 c545 (.A1(net430),
    .A2(net428),
    .A3(net439),
    .A4(net672),
    .B1(net690),
    .X(net441));
 sky130_fd_sc_hd__mux4_2 c546 (.A0(net436),
    .A1(net432),
    .A2(net907),
    .A3(net192),
    .S0(net437),
    .S1(net689),
    .X(net442));
 sky130_fd_sc_hd__a41o_1 c547 (.A1(net428),
    .A2(net442),
    .A3(net439),
    .A4(net934),
    .B1(net689),
    .X(net443));
 sky130_fd_sc_hd__mux4_1 c548 (.A0(net322),
    .A1(net427),
    .A2(net907),
    .A3(net438),
    .S0(net442),
    .S1(net672),
    .X(net444));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(net968),
    .A1(net326),
    .A2(net434),
    .A3(net442),
    .S0(net672),
    .S1(net785),
    .X(net445));
 sky130_fd_sc_hd__a41o_1 c550 (.A1(net89),
    .A2(net352),
    .A3(net76),
    .A4(net429),
    .B1(net988),
    .X(net446));
 sky130_fd_sc_hd__a41o_1 c551 (.A1(net100),
    .A2(net205),
    .A3(net446),
    .A4(net843),
    .B1(net200),
    .X(net447));
 sky130_fd_sc_hd__a41o_1 c552 (.A1(net192),
    .A2(net929),
    .A3(net334),
    .A4(net980),
    .B1(net196),
    .X(net448));
 sky130_fd_sc_hd__mux4_1 c553 (.A0(net77),
    .A1(net934),
    .A2(net950),
    .A3(net447),
    .S0(net213),
    .S1(net1014),
    .X(net449));
 sky130_fd_sc_hd__a41o_1 c554 (.A1(net427),
    .A2(net1002),
    .A3(net988),
    .A4(net698),
    .B1(net986),
    .X(net450));
 sky130_fd_sc_hd__mux4_1 c555 (.A0(net96),
    .A1(net342),
    .A2(net1003),
    .A3(net429),
    .S0(net438),
    .S1(net439),
    .X(net451));
 sky130_fd_sc_hd__sdfbbp_1 c556 (.CLK(clknet_4_8_0_clk),
    .D(net846),
    .RESET_B(net342),
    .SCD(net1009),
    .SCE(net934),
    .SET_B(net929),
    .Q(net453),
    .Q_N(net452));
 sky130_fd_sc_hd__a41o_1 c557 (.A1(net1025),
    .A2(net423),
    .A3(net209),
    .A4(net190),
    .B1(net986),
    .X(net454));
 sky130_fd_sc_hd__mux4_1 c558 (.A0(net453),
    .A1(net334),
    .A2(net703),
    .A3(net442),
    .S0(net964),
    .S1(net986),
    .X(net455));
 sky130_fd_sc_hd__mux4_2 c559 (.A0(net1022),
    .A1(net429),
    .A2(net932),
    .A3(net452),
    .S0(net934),
    .S1(net986),
    .X(net456));
 sky130_fd_sc_hd__mux4_1 c560 (.A0(net703),
    .A1(net842),
    .A2(net1053),
    .A3(net330),
    .S0(net932),
    .S1(net1068),
    .X(net457));
 sky130_fd_sc_hd__a41o_4 c561 (.A1(net95),
    .A2(net1016),
    .A3(net1015),
    .A4(net698),
    .B1(net986),
    .X(net458));
 sky130_fd_sc_hd__a41o_2 c562 (.A1(net423),
    .A2(net209),
    .A3(net1022),
    .A4(net458),
    .B1(net454),
    .X(net459));
 sky130_fd_sc_hd__a41o_1 c563 (.A1(net456),
    .A2(net339),
    .A3(net458),
    .A4(net423),
    .B1(net789),
    .X(net460));
 sky130_fd_sc_hd__a41o_2 c564 (.A1(net946),
    .A2(net944),
    .A3(net314),
    .A4(net652),
    .B1(net788),
    .X(net461));
 sky130_fd_sc_hd__sdfbbn_2 c565 (.CLK_N(clknet_4_9_0_clk),
    .D(net447),
    .RESET_B(net461),
    .SCD(net458),
    .SCE(net446),
    .SET_B(net944),
    .Q(net896),
    .Q_N(net462));
 sky130_fd_sc_hd__mux4_2 c566 (.A0(net999),
    .A1(net461),
    .A2(net213),
    .A3(net165),
    .S0(net988),
    .S1(net986),
    .X(net463));
 sky130_fd_sc_hd__a41o_1 c567 (.A1(net314),
    .A2(net462),
    .A3(net932),
    .A4(net96),
    .B1(net205),
    .X(net464));
 sky130_fd_sc_hd__sdfbbn_1 c568 (.CLK_N(clknet_4_9_0_clk),
    .D(net215),
    .RESET_B(net456),
    .SCD(net460),
    .SCE(net939),
    .SET_B(net651),
    .Q(net466),
    .Q_N(net465));
 sky130_fd_sc_hd__a41o_1 c569 (.A1(net464),
    .A2(net852),
    .A3(net466),
    .A4(net842),
    .B1(net788),
    .X(net467));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net213),
    .A1(net76),
    .A2(net454),
    .A3(net997),
    .S0(net461),
    .S1(net467),
    .X(net468));
 sky130_fd_sc_hd__mux4_1 c571 (.A0(net467),
    .A1(net429),
    .A2(net932),
    .A3(net464),
    .S0(net652),
    .S1(net790),
    .X(net469));
 sky130_fd_sc_hd__mux4_2 c572 (.A0(net375),
    .A1(net872),
    .A2(net427),
    .A3(net843),
    .S0(net684),
    .S1(net774),
    .X(net470));
 sky130_fd_sc_hd__mux4_2 c573 (.A0(net209),
    .A1(net456),
    .A2(net191),
    .A3(net458),
    .S0(net773),
    .S1(net774),
    .X(net471));
 sky130_fd_sc_hd__mux4_1 c574 (.A0(net442),
    .A1(net110),
    .A2(net345),
    .A3(net364),
    .S0(net211),
    .S1(net684),
    .X(net472));
 sky130_fd_sc_hd__mux4_1 c575 (.A0(net467),
    .A1(net873),
    .A2(net110),
    .A3(net950),
    .S0(net442),
    .S1(net773),
    .X(net473));
 sky130_fd_sc_hd__mux4_1 c576 (.A0(net342),
    .A1(net961),
    .A2(net442),
    .A3(net427),
    .S0(net338),
    .S1(net985),
    .X(net474));
 sky130_fd_sc_hd__mux4_1 c577 (.A0(net1009),
    .A1(net330),
    .A2(net460),
    .A3(net438),
    .S0(net793),
    .S1(net985),
    .X(net475));
 sky130_fd_sc_hd__mux4_2 c578 (.A0(net354),
    .A1(net459),
    .A2(net191),
    .A3(net209),
    .S0(net698),
    .S1(net793),
    .X(net476));
 sky130_fd_sc_hd__mux4_2 c579 (.A0(net863),
    .A1(net907),
    .A2(net967),
    .A3(net941),
    .S0(net944),
    .S1(net985),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c580 (.A0(net873),
    .A1(net470),
    .A2(net426),
    .A3(net364),
    .S0(net932),
    .S1(net698),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c581 (.A0(net339),
    .A1(net210),
    .A2(net330),
    .A3(net477),
    .S0(net238),
    .S1(net795),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(net869),
    .A1(net477),
    .A2(net375),
    .A3(net107),
    .S0(net684),
    .S1(net878),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c583 (.A0(net480),
    .A1(net476),
    .A2(net110),
    .A3(net98),
    .S0(net944),
    .S1(net477),
    .X(net481));
 sky130_fd_sc_hd__mux4_1 c584 (.A0(net330),
    .A1(net465),
    .A2(net375),
    .A3(net999),
    .S0(net698),
    .S1(net773),
    .X(net482));
 sky130_fd_sc_hd__mux4_1 c585 (.A0(net873),
    .A1(net364),
    .A2(net315),
    .A3(net196),
    .S0(net932),
    .S1(net793),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c586 (.A0(net454),
    .A1(net241),
    .A2(net476),
    .A3(net375),
    .S0(net828),
    .S1(clknet_1_0__leaf_net744),
    .X(net484));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(net460),
    .A1(net448),
    .A2(net364),
    .A3(net477),
    .S0(net98),
    .S1(net985),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c588 (.A0(net217),
    .A1(net869),
    .A2(net126),
    .A3(net929),
    .S0(net878),
    .S1(net793),
    .X(net486));
 sky130_fd_sc_hd__mux4_1 c589 (.A0(net983),
    .A1(net442),
    .A2(net476),
    .A3(net338),
    .S0(net895),
    .S1(net786),
    .X(net487));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(net1012),
    .A1(net426),
    .A2(net460),
    .A3(net941),
    .S0(net960),
    .S1(net985),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(net426),
    .A1(net476),
    .A2(net480),
    .A3(net324),
    .S0(net773),
    .S1(net793),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c592 (.A0(net426),
    .A1(net323),
    .A2(net477),
    .A3(net458),
    .S0(net699),
    .S1(net793),
    .X(net490));
 sky130_fd_sc_hd__mux4_2 c593 (.A0(net454),
    .A1(net490),
    .A2(net477),
    .A3(net941),
    .S0(net932),
    .S1(net686),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c594 (.A0(net205),
    .A1(net217),
    .A2(net268),
    .A3(net931),
    .S0(net989),
    .S1(net732),
    .X(net492));
 sky130_fd_sc_hd__mux4_1 c595 (.A0(net217),
    .A1(net961),
    .A2(net824),
    .A3(net891),
    .S0(net346),
    .S1(net985),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c596 (.A0(net931),
    .A1(net935),
    .A2(net427),
    .A3(net907),
    .S0(net738),
    .S1(net790),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c597 (.A0(net313),
    .A1(net959),
    .A2(net217),
    .A3(net1020),
    .S0(net735),
    .S1(clknet_1_0__leaf_net797),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c598 (.A0(net323),
    .A1(net248),
    .A2(net324),
    .A3(net714),
    .S0(net985),
    .S1(clknet_1_0__leaf_net797),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c599 (.A0(net261),
    .A1(net464),
    .A2(net313),
    .A3(net933),
    .S0(net217),
    .S1(clknet_1_0__leaf_net797),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c600 (.A0(net379),
    .A1(net1028),
    .A2(net931),
    .A3(net263),
    .S0(net239),
    .S1(net1022),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c601 (.A0(net470),
    .A1(net72),
    .A2(net315),
    .A3(net907),
    .S0(net739),
    .S1(clknet_1_0__leaf_net797),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(net196),
    .A1(net364),
    .A2(net462),
    .A3(net1017),
    .S0(net1002),
    .S1(net984),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(net268),
    .A1(net1017),
    .A2(net888),
    .A3(clknet_1_0__leaf_net495),
    .S0(net772),
    .S1(clknet_1_0__leaf_net797),
    .X(net928));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(clknet_1_1__leaf_net495),
    .A1(net843),
    .A2(net1020),
    .A3(net993),
    .S0(clknet_1_1__leaf_net710),
    .S1(net793),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net466),
    .A1(net867),
    .A2(net268),
    .A3(clknet_1_0__leaf_net495),
    .S0(net890),
    .S1(net427),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net1017),
    .A1(net458),
    .A2(clknet_1_1__leaf_net391),
    .A3(net852),
    .S0(net1003),
    .S1(net986),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(net477),
    .A1(clknet_1_0__leaf_net502),
    .A2(net915),
    .A3(net1012),
    .S0(net315),
    .S1(net772),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net863),
    .A1(net68),
    .A2(net942),
    .A3(clknet_1_1__leaf_net502),
    .S0(net737),
    .S1(clknet_1_1__leaf_net777),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c609 (.A0(clknet_1_0__leaf_net502),
    .A1(net944),
    .A2(net872),
    .A3(net346),
    .S0(net741),
    .S1(net787),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c610 (.A0(net396),
    .A1(net315),
    .A2(clknet_1_1__leaf_net502),
    .A3(net940),
    .S0(net961),
    .S1(clknet_1_1__leaf_net798),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net503),
    .A1(clknet_1_1__leaf_net502),
    .A2(clknet_1_0__leaf_net710),
    .A3(clknet_1_0__leaf_net776),
    .S0(clknet_1_0__leaf_net797),
    .S1(clknet_1_1__leaf_net798),
    .X(net508));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(net207),
    .A1(clknet_1_0__leaf_net391),
    .A2(clknet_1_1__leaf_net502),
    .A3(net989),
    .S0(net985),
    .S1(clknet_1_1__leaf_net798),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(net427),
    .A1(clknet_1_0__leaf_net502),
    .A2(net1017),
    .A3(clknet_1_0__leaf_net776),
    .S0(net787),
    .S1(clknet_1_0__leaf_net798),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(net852),
    .A1(clknet_1_1__leaf_net495),
    .A2(net347),
    .A3(net743),
    .S0(clknet_1_1__leaf_net797),
    .S1(clknet_1_0__leaf_net798),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net379),
    .A1(clknet_1_0__leaf_net511),
    .A2(net842),
    .A3(net878),
    .S0(net741),
    .S1(clknet_1_0__leaf_net798),
    .X(net512));
 sky130_fd_sc_hd__mux4_1 c616 (.A0(net199),
    .A1(net863),
    .A2(net267),
    .A3(net890),
    .S0(net728),
    .S1(clknet_1_0__leaf_net879),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(net345),
    .A1(net983),
    .A2(net413),
    .A3(net846),
    .S0(net392),
    .S1(net267),
    .X(net514));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(net324),
    .A1(net190),
    .A2(net247),
    .A3(net843),
    .S0(net1036),
    .S1(net830),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c619 (.A0(net248),
    .A1(clknet_1_0__leaf_net420),
    .A2(net956),
    .A3(net459),
    .S0(net831),
    .S1(net774),
    .X(net516));
 sky130_fd_sc_hd__mux4_2 c62 (.A0(net867),
    .A1(net858),
    .A2(net849),
    .A3(net869),
    .S0(net832),
    .S1(net865),
    .X(net0));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net68),
    .A1(net1035),
    .A2(net26),
    .A3(net949),
    .S0(net723),
    .S1(net774),
    .X(net517));
 sky130_fd_sc_hd__mux4_2 c621 (.A0(net863),
    .A1(net68),
    .A2(net835),
    .A3(net154),
    .S0(net932),
    .S1(net728),
    .X(net518));
 sky130_fd_sc_hd__mux4_2 c622 (.A0(net212),
    .A1(net16),
    .A2(net236),
    .A3(net826),
    .S0(net739),
    .S1(net756),
    .X(net519));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(net405),
    .A1(net413),
    .A2(net459),
    .A3(net82),
    .S0(net956),
    .S1(net1063),
    .X(net520));
 sky130_fd_sc_hd__mux4_2 c624 (.A0(net408),
    .A1(net956),
    .A2(net190),
    .A3(net891),
    .S0(net26),
    .S1(net987),
    .X(net521));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net843),
    .A1(net1037),
    .A2(net270),
    .A3(net931),
    .S0(net743),
    .S1(net795),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net415),
    .A1(net26),
    .A2(net518),
    .A3(net327),
    .S0(net781),
    .S1(net800),
    .X(net523));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(clknet_1_1__leaf_net420),
    .A1(net8),
    .A2(net880),
    .A3(net154),
    .S0(net742),
    .S1(net783),
    .X(net524));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net459),
    .A1(net493),
    .A2(net458),
    .A3(net69),
    .S0(net781),
    .S1(net793),
    .X(net525));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(net26),
    .A1(net518),
    .A2(net1012),
    .A3(net875),
    .S0(net678),
    .S1(net1046),
    .X(net526));
 sky130_fd_sc_hd__mux4_2 c63 (.A0(net869),
    .A1(net867),
    .A2(net859),
    .A3(net864),
    .S0(net862),
    .S1(net868),
    .X(net922));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net500),
    .A1(net846),
    .A2(net73),
    .A3(net345),
    .S0(net1014),
    .S1(net867),
    .X(net527));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net518),
    .A1(net525),
    .A2(net979),
    .A3(net997),
    .S0(net519),
    .S1(net969),
    .X(net528));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net236),
    .A1(net875),
    .A2(net471),
    .A3(net517),
    .S0(net518),
    .S1(net728),
    .X(net529));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(net471),
    .A1(net392),
    .A2(net525),
    .A3(net982),
    .S0(net740),
    .S1(net780),
    .X(net530));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net1014),
    .A1(net884),
    .A2(net728),
    .A3(net740),
    .S0(clknet_1_1__leaf_net744),
    .S1(net781),
    .X(net531));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net531),
    .A1(net896),
    .A2(net1000),
    .A3(net68),
    .S0(net889),
    .S1(net783),
    .X(net532));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net327),
    .A1(net835),
    .A2(clknet_1_1__leaf_net532),
    .A3(net519),
    .S0(net935),
    .S1(net738),
    .X(net533));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net515),
    .A1(net483),
    .A2(clknet_1_0__leaf_net532),
    .A3(net26),
    .S0(net960),
    .S1(net893),
    .X(net534));
 sky130_fd_sc_hd__mux4_2 c64 (.A0(net862),
    .A1(net860),
    .A2(net840),
    .A3(net871),
    .S0(net990),
    .S1(net858),
    .X(net1));
 sky130_fd_sc_hd__mux4_2 c65 (.A0(net832),
    .A1(net824),
    .A2(net852),
    .A3(net833),
    .S0(net995),
    .S1(net1018),
    .X(net2));
 sky130_fd_sc_hd__xnor2_1 c66 (.A(net831),
    .B(net0),
    .Y(net3));
 sky130_fd_sc_hd__a31o_1 c660 (.A1(net1005),
    .A2(net437),
    .A3(net964),
    .B1(net946),
    .X(net535));
 sky130_fd_sc_hd__a31o_1 c661 (.A1(net946),
    .A2(net80),
    .A3(net1019),
    .B1(net785),
    .X(net536));
 sky130_fd_sc_hd__a31o_1 c662 (.A1(net80),
    .A2(net437),
    .A3(net929),
    .B1(net964),
    .X(net537));
 sky130_fd_sc_hd__a41o_2 c663 (.A1(net828),
    .A2(net934),
    .A3(net929),
    .A4(net978),
    .B1(net964),
    .X(net538));
 sky130_fd_sc_hd__mux4_2 c664 (.A0(net200),
    .A1(net907),
    .A2(net437),
    .A3(net968),
    .S0(net538),
    .S1(net999),
    .X(net539));
 sky130_fd_sc_hd__a31o_1 c665 (.A1(net1004),
    .A2(net537),
    .A3(net538),
    .B1(net964),
    .X(net540));
 sky130_fd_sc_hd__a41o_2 c666 (.A1(net939),
    .A2(net978),
    .A3(net538),
    .A4(net785),
    .B1(net786),
    .X(net882));
 sky130_fd_sc_hd__a41o_1 c667 (.A1(net191),
    .A2(net1003),
    .A3(net80),
    .A4(net538),
    .B1(net1022),
    .X(net541));
 sky130_fd_sc_hd__sdfrbp_1 c668 (.CLK(clknet_4_10_0_clk),
    .D(net964),
    .RESET_B(net535),
    .SCD(net537),
    .SCE(net929),
    .Q(net543),
    .Q_N(net542));
 sky130_fd_sc_hd__a31o_1 c669 (.A1(net329),
    .A2(net535),
    .A3(net439),
    .B1(net999),
    .X(net544));
 sky130_fd_sc_hd__a21bo_1 c67 (.A1(net825),
    .A2(net1003),
    .B1_N(net1014),
    .X(net4));
 sky130_fd_sc_hd__sdfbbp_1 c670 (.CLK(clknet_4_10_0_clk),
    .D(net537),
    .RESET_B(net882),
    .SCD(net437),
    .SCE(net538),
    .SET_B(net785),
    .Q(net546),
    .Q_N(net545));
 sky130_fd_sc_hd__a31o_4 c671 (.A1(net436),
    .A2(net439),
    .A3(net978),
    .B1(net667),
    .X(net547));
 sky130_fd_sc_hd__a31o_1 c672 (.A1(net877),
    .A2(net200),
    .A3(net978),
    .B1(net667),
    .X(net548));
 sky130_fd_sc_hd__a41o_2 c673 (.A1(net68),
    .A2(net200),
    .A3(net548),
    .A4(net934),
    .B1(net439),
    .X(net549));
 sky130_fd_sc_hd__sdfbbn_1 c674 (.CLK_N(clknet_4_10_0_clk),
    .D(net535),
    .RESET_B(net548),
    .SCD(net549),
    .SCE(net964),
    .SET_B(net545),
    .Q(net551),
    .Q_N(net550));
 sky130_fd_sc_hd__a41o_1 c675 (.A1(net1005),
    .A2(net550),
    .A3(net548),
    .A4(net200),
    .B1(net667),
    .X(net552));
 sky130_fd_sc_hd__a41o_2 c676 (.A1(net552),
    .A2(net545),
    .A3(net550),
    .A4(net968),
    .B1(net547),
    .X(net553));
 sky130_fd_sc_hd__mux4_2 c677 (.A0(net548),
    .A1(net538),
    .A2(net76),
    .A3(net536),
    .S0(net542),
    .S1(net553),
    .X(net554));
 sky130_fd_sc_hd__mux4_1 c678 (.A0(net543),
    .A1(net554),
    .A2(net536),
    .A3(net316),
    .S0(net551),
    .S1(net552),
    .X(net555));
 sky130_fd_sc_hd__mux4_1 c679 (.A0(net316),
    .A1(net539),
    .A2(net552),
    .A3(net934),
    .S0(net554),
    .S1(net802),
    .X(net556));
 sky130_fd_sc_hd__xnor2_1 c68 (.A(net864),
    .B(net856),
    .Y(net5));
 sky130_fd_sc_hd__mux4_2 c680 (.A0(net551),
    .A1(net548),
    .A2(net552),
    .A3(net538),
    .S0(net667),
    .S1(net801),
    .X(net557));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(net554),
    .A1(net316),
    .A2(net557),
    .A3(net553),
    .S0(net802),
    .S1(net803),
    .X(net558));
 sky130_fd_sc_hd__mux4_1 c682 (.A0(net429),
    .A1(net552),
    .A2(net934),
    .A3(net554),
    .S0(net969),
    .S1(net1009),
    .X(net559));
 sky130_fd_sc_hd__mux4_2 c683 (.A0(net76),
    .A1(net464),
    .A2(net352),
    .A3(net831),
    .S0(net835),
    .S1(net801),
    .X(net560));
 sky130_fd_sc_hd__mux4_1 c684 (.A0(net950),
    .A1(net554),
    .A2(net352),
    .A3(net446),
    .S0(net429),
    .S1(net801),
    .X(net561));
 sky130_fd_sc_hd__mux4_1 c685 (.A0(net560),
    .A1(net538),
    .A2(net438),
    .A3(net549),
    .S0(net785),
    .S1(net1058),
    .X(net562));
 sky130_fd_sc_hd__mux4_1 c686 (.A0(net541),
    .A1(net821),
    .A2(net554),
    .A3(net786),
    .S0(net807),
    .S1(net808),
    .X(net563));
 sky130_fd_sc_hd__mux4_2 c687 (.A0(net552),
    .A1(net844),
    .A2(net934),
    .A3(net845),
    .S0(net1006),
    .S1(net808),
    .X(net564));
 sky130_fd_sc_hd__mux4_1 c688 (.A0(net98),
    .A1(net564),
    .A2(net438),
    .A3(net541),
    .S0(net993),
    .S1(net809),
    .X(net565));
 sky130_fd_sc_hd__mux4_1 c689 (.A0(net348),
    .A1(net554),
    .A2(net437),
    .A3(net994),
    .S0(net439),
    .S1(net806),
    .X(net566));
 sky130_fd_sc_hd__xnor2_4 c69 (.A(net859),
    .B(net854),
    .Y(net6));
 sky130_fd_sc_hd__mux4_2 c690 (.A0(net934),
    .A1(net542),
    .A2(net547),
    .A3(net830),
    .S0(net786),
    .S1(net792),
    .X(net567));
 sky130_fd_sc_hd__mux4_1 c691 (.A0(net216),
    .A1(net1019),
    .A2(net788),
    .A3(net805),
    .S0(net806),
    .S1(net808),
    .X(net568));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(net329),
    .A1(net541),
    .A2(net461),
    .A3(net939),
    .S0(net554),
    .S1(net1051),
    .X(net569));
 sky130_fd_sc_hd__mux4_1 c693 (.A0(net819),
    .A1(net568),
    .A2(net554),
    .A3(net830),
    .S0(net80),
    .S1(net681),
    .X(net570));
 sky130_fd_sc_hd__mux4_2 c694 (.A0(net352),
    .A1(net845),
    .A2(net348),
    .A3(net441),
    .S0(net429),
    .S1(net808),
    .X(net571));
 sky130_fd_sc_hd__mux4_2 c695 (.A0(net543),
    .A1(net329),
    .A2(net107),
    .A3(net571),
    .S0(net694),
    .S1(net801),
    .X(net883));
 sky130_fd_sc_hd__mux4_2 c696 (.A0(net334),
    .A1(net946),
    .A2(net1005),
    .A3(net978),
    .S0(net845),
    .S1(net805),
    .X(net572));
 sky130_fd_sc_hd__mux4_1 c697 (.A0(net446),
    .A1(net841),
    .A2(net557),
    .A3(net883),
    .S0(net694),
    .S1(net1064),
    .X(net573));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(net553),
    .A1(net883),
    .A2(net978),
    .A3(net681),
    .S0(net809),
    .S1(net812),
    .X(net574));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(net461),
    .A1(net571),
    .A2(net536),
    .A3(net568),
    .S0(net553),
    .S1(net805),
    .X(net575));
 sky130_fd_sc_hd__a21bo_1 c70 (.A1(net997),
    .A2(net4),
    .B1_N(net859),
    .X(net7));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net224),
    .A1(net883),
    .A2(net76),
    .A3(net554),
    .S0(net813),
    .S1(net814),
    .X(net576));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(net536),
    .A1(net571),
    .A2(clknet_1_0__leaf_net711),
    .A3(net791),
    .S0(net806),
    .S1(net814),
    .X(net577));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net572),
    .A1(clknet_1_0__leaf_net577),
    .A2(net553),
    .A3(net883),
    .S0(net698),
    .S1(net814),
    .X(net578));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(clknet_1_0__leaf_net577),
    .A1(net541),
    .A2(net693),
    .A3(net810),
    .S0(net814),
    .S1(net815),
    .X(net579));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net820),
    .A1(net242),
    .A2(net567),
    .A3(net572),
    .S0(net950),
    .S1(net681),
    .X(net580));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(net867),
    .A1(net939),
    .A2(net693),
    .A3(net986),
    .S0(clknet_1_0__leaf_net796),
    .S1(net801),
    .X(net581));
 sky130_fd_sc_hd__mux4_1 c706 (.A0(net538),
    .A1(net1004),
    .A2(net936),
    .A3(net947),
    .S0(net883),
    .S1(net458),
    .X(net582));
 sky130_fd_sc_hd__mux4_2 c707 (.A0(net98),
    .A1(net107),
    .A2(net247),
    .A3(net786),
    .S0(net794),
    .S1(net807),
    .X(net583));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(net996),
    .A1(net965),
    .A2(net107),
    .A3(net547),
    .S0(net768),
    .S1(net804),
    .X(net584));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(net98),
    .A1(net437),
    .A2(net463),
    .A3(net1006),
    .S0(clknet_1_0__leaf_net711),
    .S1(net986),
    .X(net585));
 sky130_fd_sc_hd__xnor2_4 c71 (.A(net821),
    .B(net1017),
    .Y(net8));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net0),
    .A1(net1013),
    .A2(net547),
    .A3(net583),
    .S0(net126),
    .S1(clknet_1_0__leaf_net744),
    .X(net586));
 sky130_fd_sc_hd__mux4_2 c711 (.A0(net110),
    .A1(net491),
    .A2(net584),
    .A3(net242),
    .S0(net962),
    .S1(net437),
    .X(net587));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net557),
    .A1(net110),
    .A2(net448),
    .A3(net126),
    .S0(net191),
    .S1(net807),
    .X(net588));
 sky130_fd_sc_hd__mux4_1 c713 (.A0(net572),
    .A1(net491),
    .A2(net587),
    .A3(net895),
    .S0(net750),
    .S1(net768),
    .X(net589));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(net338),
    .A1(net241),
    .A2(net882),
    .A3(net978),
    .S0(clknet_1_1__leaf_net577),
    .S1(net804),
    .X(net590));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net437),
    .A1(net1013),
    .A2(net98),
    .A3(net822),
    .S0(net567),
    .S1(net816),
    .X(net591));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net587),
    .A1(net824),
    .A2(net463),
    .A3(net583),
    .S0(net564),
    .S1(net772),
    .X(net592));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net571),
    .A1(net567),
    .A2(net587),
    .A3(net819),
    .S0(net786),
    .S1(net788),
    .X(net593));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(net126),
    .A1(net587),
    .A2(net968),
    .A3(net786),
    .S0(clknet_1_1__leaf_net796),
    .S1(net816),
    .X(net594));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net1006),
    .A1(net845),
    .A2(net239),
    .A3(net572),
    .S0(net107),
    .S1(clknet_1_0__leaf_net775),
    .X(net595));
 sky130_fd_sc_hd__a21bo_4 c72 (.A1(net0),
    .A2(net860),
    .B1_N(net1),
    .X(net9));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net585),
    .A1(net347),
    .A2(net0),
    .A3(net491),
    .S0(net786),
    .S1(clknet_1_0__leaf_net817),
    .X(net596));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net448),
    .A1(net580),
    .A2(net347),
    .A3(net583),
    .S0(net587),
    .S1(net806),
    .X(net597));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net567),
    .A1(net338),
    .A2(net557),
    .A3(net978),
    .S1(net746),
    .X(net598));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net72),
    .A1(net587),
    .A2(net1070),
    .A3(net1066),
    .S0(net807),
    .S1(net1047),
    .X(net599));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net491),
    .A1(net895),
    .A2(net747),
    .A3(net750),
    .S0(net815),
    .S1(clknet_1_0__leaf_net817),
    .X(net600));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net241),
    .A1(net546),
    .A2(net220),
    .A3(clknet_1_0__leaf_net600),
    .S0(net715),
    .S1(net813),
    .X(net601));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net15),
    .A1(net966),
    .A2(net0),
    .A3(net750),
    .S0(clknet_1_1__leaf_net797),
    .S1(net802),
    .X(net602));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(clknet_1_1__leaf_net577),
    .A1(net931),
    .A2(net219),
    .A3(net560),
    .S0(net882),
    .S1(net686),
    .X(net603));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net591),
    .A1(net581),
    .A2(net549),
    .A3(net845),
    .S0(net720),
    .S1(net806),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(net490),
    .A1(net960),
    .A2(net584),
    .A3(net935),
    .S0(clknet_1_0__leaf_net775),
    .S1(clknet_1_0__leaf_net818),
    .X(net605));
 sky130_fd_sc_hd__xnor2_4 c73 (.A(net834),
    .B(net864),
    .Y(net10));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net841),
    .A1(net501),
    .A2(net211),
    .A3(net933),
    .S0(net947),
    .S1(net739),
    .X(net606));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net497),
    .A1(net984),
    .A2(net857),
    .A3(net458),
    .S0(clknet_1_0__leaf_net602),
    .S1(net539),
    .X(net607));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(net549),
    .A1(net547),
    .A2(net736),
    .A3(net746),
    .S0(net985),
    .S1(clknet_1_1__leaf_net817),
    .X(net608));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net824),
    .A1(net848),
    .A2(net512),
    .A3(net883),
    .S0(net821),
    .S1(net463),
    .X(net609));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(clknet_1_1__leaf_net398),
    .A1(net989),
    .A2(clknet_1_1__leaf_net710),
    .A3(net716),
    .S0(net736),
    .S1(net802),
    .X(net610));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net936),
    .A1(net933),
    .A2(net326),
    .A3(net88),
    .S0(clknet_1_1__leaf_net711),
    .S1(net985),
    .X(net611));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(net347),
    .A1(net219),
    .A2(net564),
    .A3(net936),
    .S0(clknet_1_0__leaf_net600),
    .S1(net743),
    .X(net612));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net463),
    .A1(clknet_1_0__leaf_net511),
    .A2(net539),
    .A3(net828),
    .S0(net989),
    .S1(clknet_1_1__leaf_net797),
    .X(net613));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net239),
    .A1(net959),
    .A2(net915),
    .A3(net591),
    .S0(net269),
    .S1(net772),
    .X(net614));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(net326),
    .A1(net936),
    .A2(clknet_1_1__leaf_net879),
    .A3(clknet_1_1__leaf_net776),
    .S0(net810),
    .S1(clknet_1_0__leaf_net818),
    .X(net615));
 sky130_fd_sc_hd__xnor2_2 c74 (.A(net7),
    .B(net858),
    .Y(net11));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(net583),
    .A1(net831),
    .A2(net857),
    .A3(net959),
    .S0(net720),
    .S1(net802),
    .X(net616));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(net606),
    .A1(net560),
    .A2(net933),
    .A3(net966),
    .S0(net929),
    .S1(clknet_1_1__leaf_net797),
    .X(net617));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(net546),
    .A1(net857),
    .A2(net931),
    .A3(net583),
    .S0(net886),
    .S1(net806),
    .X(net618));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(clknet_1_0__leaf_net611),
    .A1(clknet_1_1__leaf_net600),
    .A2(clknet_1_0__leaf_net610),
    .A3(net915),
    .S0(clknet_1_0__leaf_net775),
    .S1(clknet_1_0__leaf_net818),
    .X(net619));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(clknet_1_1__leaf_net611),
    .A1(net979),
    .A2(clknet_1_1__leaf_net595),
    .A3(net720),
    .S0(net886),
    .S1(net739),
    .X(net887));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(clknet_1_0__leaf_net615),
    .A1(net0),
    .A2(net583),
    .A3(net845),
    .S0(clknet_1_0__leaf_net879),
    .S1(net806),
    .X(net620));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net549),
    .A1(clknet_1_1__leaf_net615),
    .A2(clknet_1_1__leaf_net511),
    .A3(net716),
    .S0(net720),
    .S1(net738),
    .X(net621));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(net564),
    .A1(net621),
    .A2(net219),
    .A3(net105),
    .S0(net685),
    .S1(net806),
    .X(net622));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net959),
    .A1(net861),
    .A2(net392),
    .A3(net877),
    .S0(net1001),
    .S1(net844),
    .X(net623));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net458),
    .A1(net623),
    .A2(net1023),
    .A3(net935),
    .S0(clknet_1_1__leaf_net711),
    .S1(net715),
    .X(net624));
 sky130_fd_sc_hd__a21bo_2 c75 (.A1(net823),
    .A2(net870),
    .B1_N(net852),
    .X(net12));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(net539),
    .A1(net267),
    .A2(net839),
    .A3(net624),
    .S0(net1041),
    .S1(clknet_1_1__leaf_net818),
    .X(net625));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(clknet_1_0__leaf_net595),
    .A1(net831),
    .A2(net513),
    .A3(clknet_1_1__leaf_net608),
    .S0(net521),
    .S1(clknet_1_1__leaf_net775),
    .X(net626));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net263),
    .A1(net211),
    .A2(net969),
    .A3(net69),
    .S0(net122),
    .S1(net737),
    .X(net627));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(clknet_1_1__leaf_net602),
    .A1(net1028),
    .A2(net1020),
    .A3(clknet_1_0__leaf_net608),
    .S0(net893),
    .S1(net811),
    .X(net628));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net269),
    .A1(net993),
    .A2(net861),
    .A3(net932),
    .S0(net211),
    .S1(net736),
    .X(net629));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net1001),
    .A1(net628),
    .A2(net881),
    .A3(net1037),
    .S0(net737),
    .S1(net756),
    .X(net630));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net932),
    .A1(net940),
    .A2(net909),
    .A3(net979),
    .S0(net722),
    .S1(net743),
    .X(net631));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(clknet_1_1__leaf_net610),
    .A1(net627),
    .A2(net418),
    .A3(net883),
    .S0(clknet_1_1__leaf_net775),
    .S1(net811),
    .X(net632));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net839),
    .A1(net906),
    .A2(net886),
    .A3(net893),
    .S0(net793),
    .S1(net815),
    .X(net633));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net82),
    .A1(net633),
    .A2(net8),
    .A3(net828),
    .S0(net761),
    .S1(clknet_1_1__leaf_net818),
    .X(net634));
 sky130_fd_sc_hd__a21bo_4 c76 (.A1(net9),
    .A2(net1011),
    .B1_N(net6),
    .X(net13));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net418),
    .A1(net15),
    .A2(net392),
    .A3(net450),
    .S0(net737),
    .S1(net987),
    .X(net635));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net635),
    .A1(net867),
    .A2(net527),
    .A3(net634),
    .S0(net968),
    .S1(net940),
    .X(net636));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net247),
    .A1(net884),
    .A2(net907),
    .A3(net736),
    .S0(net740),
    .S1(net750),
    .X(net637));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(net317),
    .A1(net122),
    .A2(net16),
    .A3(net521),
    .S0(net247),
    .S1(net915),
    .X(net638));
 sky130_fd_sc_hd__mux4_1 c764 (.A0(net400),
    .A1(net979),
    .A2(net605),
    .A3(net68),
    .S0(net15),
    .S1(net966),
    .X(net639));
 sky130_fd_sc_hd__mux4_1 c765 (.A0(net270),
    .A1(net8),
    .A2(clknet_1_1__leaf_net398),
    .A3(net638),
    .S0(clknet_1_0__leaf_net595),
    .S1(net740),
    .X(net640));
 sky130_fd_sc_hd__mux4_1 c766 (.A0(net88),
    .A1(net1041),
    .A2(net622),
    .A3(net637),
    .S0(net959),
    .S1(net861),
    .X(net641));
 sky130_fd_sc_hd__mux4_1 c767 (.A0(net517),
    .A1(net839),
    .A2(clknet_1_1__leaf_net398),
    .A3(net695),
    .S0(net704),
    .S1(net738),
    .X(net642));
 sky130_fd_sc_hd__mux4_1 c768 (.A0(net547),
    .A1(net1020),
    .A2(net519),
    .A3(net639),
    .S0(net642),
    .S1(net742),
    .X(net643));
 sky130_fd_sc_hd__mux4_1 c769 (.A0(net1020),
    .A1(net638),
    .A2(net678),
    .A3(net722),
    .S0(net781),
    .S1(net793),
    .X(net644));
 sky130_fd_sc_hd__xnor2_2 c77 (.A(net827),
    .B(net10),
    .Y(net14));
 sky130_fd_sc_hd__a21bo_2 c78 (.A1(net10),
    .A2(net3),
    .B1_N(net9),
    .X(net15));
 sky130_fd_sc_hd__a21bo_2 c79 (.A1(net15),
    .A2(net12),
    .B1_N(net875),
    .X(net16));
 sky130_fd_sc_hd__a21bo_1 c80 (.A1(net13),
    .A2(net6),
    .B1_N(net866),
    .X(net17));
 sky130_fd_sc_hd__a31o_4 c81 (.A1(net14),
    .A2(net871),
    .A3(net11),
    .B1(net970),
    .X(net18));
 sky130_fd_sc_hd__mux4_2 c82 (.A0(net12),
    .A1(net18),
    .A2(net852),
    .A3(net864),
    .S0(net10),
    .S1(net970),
    .X(net19));
 sky130_fd_sc_hd__a41o_4 c83 (.A1(net16),
    .A2(net18),
    .A3(net970),
    .A4(net13),
    .B1(net19),
    .X(net20));
 sky130_fd_sc_hd__mux4_2 c84 (.A0(net20),
    .A1(net856),
    .A2(net970),
    .A3(net8),
    .S0(net12),
    .S1(net857),
    .X(net21));
 sky130_fd_sc_hd__mux4_2 c85 (.A0(net19),
    .A1(net5),
    .A2(net12),
    .A3(net13),
    .S0(net859),
    .S1(net21),
    .X(net22));
 sky130_fd_sc_hd__a31o_4 c86 (.A1(net6),
    .A2(net951),
    .A3(net8),
    .B1(net970),
    .X(net23));
 sky130_fd_sc_hd__mux4_2 c87 (.A0(net973),
    .A1(net3),
    .A2(net23),
    .A3(net951),
    .S0(net4),
    .S1(net21),
    .X(net24));
 sky130_fd_sc_hd__a21bo_4 c88 (.A1(net850),
    .A2(net13),
    .B1_N(net24),
    .X(net25));
 sky130_fd_sc_hd__a21bo_4 c89 (.A1(net1011),
    .A2(net866),
    .B1_N(net972),
    .X(net26));
 sky130_fd_sc_hd__a21bo_1 c90 (.A1(net874),
    .A2(net858),
    .B1_N(net1014),
    .X(net27));
 sky130_fd_sc_hd__a31o_1 c91 (.A1(net838),
    .A2(net854),
    .A3(net18),
    .B1(net1007),
    .X(net28));
 sky130_fd_sc_hd__a31o_2 c92 (.A1(net3),
    .A2(net1014),
    .A3(net28),
    .B1(net837),
    .X(net29));
 sky130_fd_sc_hd__a21bo_2 c93 (.A1(net7),
    .A2(net1021),
    .B1_N(net973),
    .X(net30));
 sky130_fd_sc_hd__a21bo_4 c94 (.A1(net843),
    .A2(net2),
    .B1_N(net862),
    .X(net31));
 sky130_fd_sc_hd__a21bo_1 c95 (.A1(net13),
    .A2(net867),
    .B1_N(net24),
    .X(net32));
 sky130_fd_sc_hd__a21bo_1 c96 (.A1(net12),
    .A2(net30),
    .B1_N(net867),
    .X(net33));
 sky130_fd_sc_hd__a21bo_1 c97 (.A1(net1018),
    .A2(net857),
    .B1_N(net26),
    .X(net34));
 sky130_fd_sc_hd__a21bo_2 c98 (.A1(net866),
    .A2(net11),
    .B1_N(net12),
    .X(net35));
 sky130_fd_sc_hd__a21bo_4 c99 (.A1(net4),
    .A2(net25),
    .B1_N(net856),
    .X(net36));
 sky130_fd_sc_hd__a41o_1 merge790 (.A1(net333),
    .A2(net221),
    .A3(net206),
    .A4(net336),
    .B1(net337),
    .X(net645));
 sky130_fd_sc_hd__mux4_1 merge791 (.A0(net331),
    .A1(net318),
    .A2(net314),
    .A3(net207),
    .S0(net431),
    .S1(net999),
    .X(net646));
 sky130_fd_sc_hd__xnor2_1 merge792 (.A(net401),
    .B(net411),
    .Y(net647));
 sky130_fd_sc_hd__xnor2_1 merge793 (.A(net380),
    .B(net381),
    .Y(net648));
 sky130_fd_sc_hd__xnor2_1 merge794 (.A(net230),
    .B(net226),
    .Y(net649));
 sky130_fd_sc_hd__xnor2_1 merge795 (.A(net294),
    .B(net296),
    .Y(net650));
 sky130_fd_sc_hd__dfrbp_1 merge796 (.CLK(clknet_4_10_0_clk),
    .D(net468),
    .RESET_B(net457),
    .Q(net652),
    .Q_N(net651));
 sky130_fd_sc_hd__xnor2_1 merge797 (.A(net604),
    .B(net607),
    .Y(net653));
 sky130_fd_sc_hd__dfrbp_1 merge798 (.CLK(clknet_4_9_0_clk),
    .D(net357),
    .RESET_B(net372),
    .Q(net655),
    .Q_N(net654));
 sky130_fd_sc_hd__xnor2_1 merge799 (.A(net484),
    .B(net485),
    .Y(net656));
 sky130_fd_sc_hd__xnor2_1 merge800 (.A(net272),
    .B(net252),
    .Y(net657));
 sky130_fd_sc_hd__xnor2_1 merge801 (.A(net250),
    .B(net243),
    .Y(net658));
 sky130_fd_sc_hd__xnor2_1 merge802 (.A(net592),
    .B(net593),
    .Y(net659));
 sky130_fd_sc_hd__xnor2_1 merge803 (.A(net644),
    .B(net625),
    .Y(net660));
 sky130_fd_sc_hd__xnor2_1 merge804 (.A(net514),
    .B(net520),
    .Y(net661));
 sky130_fd_sc_hd__xnor2_1 merge805 (.A(net286),
    .B(net283),
    .Y(net662));
 sky130_fd_sc_hd__dfrtn_1 merge806 (.CLK_N(clknet_4_8_0_clk),
    .D(net645),
    .RESET_B(net349),
    .Q(net663));
 sky130_fd_sc_hd__dfrtp_4 merge807 (.CLK(clknet_4_3_0_clk),
    .D(net148),
    .RESET_B(net146),
    .Q(net664));
 sky130_fd_sc_hd__xnor2_1 merge808 (.A(net64),
    .B(net63),
    .Y(net665));
 sky130_fd_sc_hd__xnor2_1 merge809 (.A(net159),
    .B(net163),
    .Y(net666));
 sky130_fd_sc_hd__dfrtp_2 merge810 (.CLK(clknet_4_10_0_clk),
    .D(net540),
    .RESET_B(net544),
    .Q(net667));
 sky130_fd_sc_hd__xnor2_1 merge811 (.A(net183),
    .B(net188),
    .Y(net668));
 sky130_fd_sc_hd__xnor2_1 merge812 (.A(net566),
    .B(net578),
    .Y(net669));
 sky130_fd_sc_hd__xnor2_1 merge813 (.A(net421),
    .B(net422),
    .Y(net670));
 sky130_fd_sc_hd__xnor2_1 merge814 (.A(net492),
    .B(net498),
    .Y(net671));
 sky130_fd_sc_hd__dfrtp_1 merge815 (.CLK(clknet_4_8_0_clk),
    .D(net424),
    .RESET_B(net443),
    .Q(net672));
 sky130_fd_sc_hd__xnor2_1 merge816 (.A(net416),
    .B(net311),
    .Y(net673));
 sky130_fd_sc_hd__dfsbp_2 merge817 (.CLK(clknet_4_5_0_clk),
    .SET_B(net666),
    .Q(net675),
    .Q_N(net674));
 sky130_fd_sc_hd__dfsbp_2 merge818 (.CLK(clknet_4_3_0_clk),
    .D(net255),
    .SET_B(net229),
    .Q(net677),
    .Q_N(net676));
 sky130_fd_sc_hd__dfstp_1 merge819 (.CLK(clknet_4_13_0_clk),
    .D(net524),
    .SET_B(net643),
    .Q(net678));
 sky130_fd_sc_hd__xnor2_1 merge820 (.A(net522),
    .B(net309),
    .Y(net679));
 sky130_fd_sc_hd__xnor2_1 merge821 (.A(net303),
    .B(net298),
    .Y(net680));
 sky130_fd_sc_hd__dfstp_1 merge822 (.CLK(clknet_4_11_0_clk),
    .D(net579),
    .SET_B(net569),
    .Q(net681));
 sky130_fd_sc_hd__xnor2_1 merge823 (.A(net487),
    .B(net620),
    .Y(net682));
 sky130_fd_sc_hd__xnor2_1 merge824 (.A(net488),
    .B(net619),
    .Y(net683));
 sky130_fd_sc_hd__dfstp_2 merge825 (.CLK(clknet_4_2_0_clk),
    .D(net244),
    .SET_B(net370),
    .Q(net684));
 sky130_fd_sc_hd__dlrbn_1 merge826 (.D(net489),
    .GATE_N(clknet_4_14_0_clk),
    .RESET_B(net683),
    .Q(net686),
    .Q_N(net685));
 sky130_fd_sc_hd__xnor2_1 merge827 (.A(net660),
    .B(net507),
    .Y(net687));
 sky130_fd_sc_hd__xnor2_1 merge828 (.A(net523),
    .B(net641),
    .Y(net688));
 sky130_fd_sc_hd__dlrbn_1 merge829 (.D(net646),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net440),
    .Q(net690),
    .Q_N(net689));
 sky130_fd_sc_hd__dlrbp_1 merge830 (.D(net662),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net290),
    .Q(net692),
    .Q_N(net691));
 sky130_fd_sc_hd__dlrbp_1 merge831 (.D(net565),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net669),
    .Q(net694),
    .Q_N(net693));
 sky130_fd_sc_hd__dlrtn_1 merge832 (.D(net673),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net647),
    .Q(net908));
 sky130_fd_sc_hd__dlrtn_1 merge833 (.D(net147),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net143),
    .Q(net695));
 sky130_fd_sc_hd__xnor2_1 merge834 (.A(net305),
    .B(net680),
    .Y(net696));
 sky130_fd_sc_hd__dlrtn_2 merge835 (.D(net649),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net228),
    .Q(net697));
 sky130_fd_sc_hd__dlrtp_4 merge836 (.D(net344),
    .GATE(clknet_4_9_0_clk),
    .RESET_B(net351),
    .Q(net698));
 sky130_fd_sc_hd__dlrtp_2 merge837 (.D(net237),
    .GATE(clknet_4_2_0_clk),
    .RESET_B(net245),
    .Q(net699));
 sky130_fd_sc_hd__xnor2_1 merge838 (.A(net504),
    .B(net528),
    .Y(net700));
 sky130_fd_sc_hd__xnor2_1 merge839 (.A(net529),
    .B(net640),
    .Y(net701));
 sky130_fd_sc_hd__dlrtp_1 merge840 (.D(net668),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net182),
    .Q(net702));
 sky130_fd_sc_hd__edfxbp_1 merge841 (.CLK(clknet_4_14_0_clk),
    .DE(net659),
    .Q(net704),
    .Q_N(net598));
 sky130_fd_sc_hd__xnor2_1 merge842 (.A(net530),
    .B(net636),
    .Y(net705));
 sky130_fd_sc_hd__edfxtp_1 merge843 (.CLK(clknet_4_4_0_clk),
    .D(net665),
    .DE(net650),
    .Q(net927));
 sky130_fd_sc_hd__xnor2_1 merge844 (.A(net533),
    .B(net534),
    .Y(net706));
 sky130_fd_sc_hd__xnor2_1 merge845 (.A(net499),
    .B(net510),
    .Y(net707));
 sky130_fd_sc_hd__xnor2_1 merge846 (.A(net508),
    .B(net505),
    .Y(net708));
 sky130_fd_sc_hd__sdlclkp_1 merge847 (.CLK(clknet_4_0_0_clk),
    .GATE(net175),
    .GCLK(net709));
 sky130_fd_sc_hd__sdlclkp_2 merge848 (.CLK(clknet_4_6_0_clk),
    .GATE(net397),
    .SCE(net383),
    .GCLK(net710));
 sky130_fd_sc_hd__sdlclkp_4 merge849 (.CLK(clknet_4_11_0_clk),
    .GATE(net574),
    .SCE(net601),
    .GCLK(net711));
 sky130_fd_sc_hd__xnor2_1 merge850 (.A(net509),
    .B(net632),
    .Y(net712));
 sky130_fd_sc_hd__dfrbp_1 merge851 (.CLK(clknet_4_6_0_clk),
    .D(net256),
    .RESET_B(net282),
    .Q(net714),
    .Q_N(net713));
 sky130_fd_sc_hd__dfrbp_2 merge852 (.CLK(clknet_4_14_0_clk),
    .D(net481),
    .RESET_B(net599),
    .Q(net716),
    .Q_N(net715));
 sky130_fd_sc_hd__xnor2_1 merge853 (.A(net618),
    .B(net609),
    .Y(net717));
 sky130_fd_sc_hd__xnor2_1 merge854 (.A(net617),
    .B(net612),
    .Y(net718));
 sky130_fd_sc_hd__xnor2_1 merge855 (.A(net613),
    .B(net616),
    .Y(net719));
 sky130_fd_sc_hd__dfrtn_1 merge856 (.CLK_N(clknet_4_15_0_clk),
    .D(net582),
    .RESET_B(net718),
    .Q(net720));
 sky130_fd_sc_hd__dfrtp_4 merge857 (.CLK(clknet_4_0_0_clk),
    .D(net260),
    .RESET_B(net181),
    .Q(net899));
 sky130_fd_sc_hd__dfrtp_2 merge858 (.CLK(clknet_4_14_0_clk),
    .D(net474),
    .RESET_B(net712),
    .Q(net878));
 sky130_fd_sc_hd__dfrtp_1 merge859 (.CLK(clknet_4_0_0_clk),
    .D(net249),
    .Q(net251));
 sky130_fd_sc_hd__dfsbp_1 merge860 (.CLK(clknet_4_6_0_clk),
    .D(net409),
    .SET_B(net706),
    .Q(net723),
    .Q_N(net722));
 sky130_fd_sc_hd__dfsbp_1 merge861 (.CLK(clknet_4_6_0_clk),
    .D(net412),
    .SET_B(net410),
    .Q(net725),
    .Q_N(net724));
 sky130_fd_sc_hd__dfstp_1 merge862 (.CLK(clknet_4_15_0_clk),
    .D(net719),
    .SET_B(net717),
    .Q(net886));
 sky130_fd_sc_hd__xnor2_1 merge863 (.A(net631),
    .B(net626),
    .Y(net726));
 sky130_fd_sc_hd__dfstp_2 merge864 (.CLK(clknet_4_0_0_clk),
    .D(net658),
    .SET_B(net356),
    .Q(net727));
 sky130_fd_sc_hd__dfstp_1 merge865 (.CLK(clknet_4_7_0_clk),
    .D(net402),
    .SET_B(net399),
    .Q(net728));
 sky130_fd_sc_hd__dlrbn_1 merge866 (.D(net362),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net648),
    .Q(net730),
    .Q_N(net729));
 sky130_fd_sc_hd__dlrbn_1 merge867 (.D(net265),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net273),
    .Q(net732),
    .Q_N(net731));
 sky130_fd_sc_hd__xnor2_1 merge868 (.A(net630),
    .B(net629),
    .Y(net733));
 sky130_fd_sc_hd__dlrbp_1 merge869 (.D(net670),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net277),
    .Q(net930),
    .Q_N(net734));
 sky130_fd_sc_hd__dlrbp_2 merge870 (.D(net657),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net696),
    .Q(net735),
    .Q_N(net897));
 sky130_fd_sc_hd__dlrtn_1 merge871 (.D(net590),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net726),
    .Q(net736));
 sky130_fd_sc_hd__dlrtn_1 merge872 (.D(net671),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net733),
    .Q(net737));
 sky130_fd_sc_hd__dlrtn_2 merge873 (.D(net682),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net701),
    .Q(net738));
 sky130_fd_sc_hd__dlrtp_2 merge874 (.D(net496),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net653),
    .Q(net739));
 sky130_fd_sc_hd__dlrtp_1 merge875 (.D(net656),
    .GATE(clknet_4_12_0_clk),
    .RESET_B(net486),
    .Q(net895));
 sky130_fd_sc_hd__dlrtp_1 merge876 (.D(net705),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net700),
    .Q(net740));
 sky130_fd_sc_hd__edfxbp_1 merge877 (.CLK(clknet_4_13_0_clk),
    .D(net688),
    .DE(net707),
    .Q(net742),
    .Q_N(net741));
 sky130_fd_sc_hd__edfxtp_1 merge878 (.CLK(clknet_4_13_0_clk),
    .D(net687),
    .DE(net708),
    .Q(net743));
 sky130_fd_sc_hd__sdlclkp_1 merge879 (.CLK(clknet_4_15_0_clk),
    .GATE(net479),
    .SCE(net614),
    .GCLK(net879));
 sky130_fd_sc_hd__sdlclkp_2 merge880 (.CLK(clknet_4_12_0_clk),
    .GATE(net679),
    .SCE(net482),
    .GCLK(net744));
 sky130_fd_sc_hd__sdlclkp_4 merge881 (.CLK(clknet_4_0_0_clk),
    .GATE(net234),
    .GCLK(net235));
 sky130_fd_sc_hd__dfrbp_1 merge882 (.CLK(clknet_4_14_0_clk),
    .D(net597),
    .RESET_B(net596),
    .Q(net747),
    .Q_N(net746));
 sky130_fd_sc_hd__dfrbp_2 merge883 (.CLK(clknet_4_4_0_clk),
    .D(net184),
    .RESET_B(net295),
    .Q(net749),
    .Q_N(net748));
 sky130_fd_sc_hd__dfrtn_1 merge884 (.CLK_N(clknet_4_13_0_clk),
    .D(net661),
    .RESET_B(net526),
    .Q(net893));
 sky130_fd_sc_hd__dfrtp_2 merge885 (.CLK(clknet_4_14_0_clk),
    .D(net588),
    .RESET_B(net586),
    .Q(net750));
 sky130_fd_sc_hd__dfxbp_1 s886 (.CLK(clknet_4_1_0_clk),
    .D(net57),
    .Q(net752),
    .Q_N(net751));
 sky130_fd_sc_hd__dfxbp_1 s887 (.CLK(clknet_4_1_0_clk),
    .D(net144),
    .Q(net754),
    .Q_N(net753));
 sky130_fd_sc_hd__dfxtp_1 s888 (.CLK(clknet_4_4_0_clk),
    .D(net153),
    .Q(net755));
 sky130_fd_sc_hd__dfxtp_2 s889 (.CLK(clknet_4_5_0_clk),
    .D(net167),
    .Q(net756));
 sky130_fd_sc_hd__dfxtp_2 s890 (.CLK(clknet_4_5_0_clk),
    .D(net168),
    .Q(net757));
 sky130_fd_sc_hd__dlclkp_1 s891 (.CLK(clknet_4_5_0_clk),
    .GATE(net169),
    .GCLK(net758));
 sky130_fd_sc_hd__dlclkp_2 s892 (.CLK(clknet_4_0_0_clk),
    .GATE(net172),
    .GCLK(net759));
 sky130_fd_sc_hd__dlclkp_4 s893 (.CLK(clknet_4_0_0_clk),
    .GATE(net178),
    .GCLK(net901));
 sky130_fd_sc_hd__dlxbn_2 s894 (.D(net253),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net761),
    .Q_N(net760));
 sky130_fd_sc_hd__dlxbn_1 s895 (.D(net274),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net920),
    .Q_N(net762));
 sky130_fd_sc_hd__dlxbp_1 s896 (.D(net287),
    .GATE(clknet_4_7_0_clk),
    .Q(net925),
    .Q_N(net763));
 sky130_fd_sc_hd__dlxtn_1 s897 (.D(net288),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net764));
 sky130_fd_sc_hd__dlxtn_1 s898 (.D(net291),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net765));
 sky130_fd_sc_hd__dlxtn_1 s899 (.D(net301),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net766));
 sky130_fd_sc_hd__dlxtp_1 s900 (.D(net332),
    .GATE(clknet_4_8_0_clk),
    .Q(net767));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s901 (.D(net361),
    .SLEEP_B(clknet_4_9_0_clk),
    .Q(net768));
 sky130_fd_sc_hd__dfxbp_1 s902 (.CLK(clknet_4_9_0_clk),
    .D(net363),
    .Q(net770),
    .Q_N(net769));
 sky130_fd_sc_hd__dfxbp_1 s903 (.CLK(clknet_4_6_0_clk),
    .D(net366),
    .Q(net921),
    .Q_N(net771));
 sky130_fd_sc_hd__dfxtp_2 s904 (.CLK(clknet_4_3_0_clk),
    .D(net369),
    .Q(net772));
 sky130_fd_sc_hd__dfxtp_2 s905 (.CLK(clknet_4_12_0_clk),
    .D(net373),
    .Q(net773));
 sky130_fd_sc_hd__dfxtp_2 s906 (.CLK(clknet_4_12_0_clk),
    .D(net374),
    .Q(net774));
 sky130_fd_sc_hd__dlclkp_1 s907 (.CLK(clknet_4_12_0_clk),
    .GATE(net376),
    .GCLK(net775));
 sky130_fd_sc_hd__dlclkp_2 s908 (.CLK(clknet_4_12_0_clk),
    .GATE(net385),
    .GCLK(net776));
 sky130_fd_sc_hd__dlclkp_4 s909 (.CLK(clknet_4_13_0_clk),
    .GATE(net388),
    .GCLK(net777));
 sky130_fd_sc_hd__dlxbn_1 s910 (.D(net394),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net779),
    .Q_N(net778));
 sky130_fd_sc_hd__dlxbn_1 s911 (.D(net404),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net781),
    .Q_N(net780));
 sky130_fd_sc_hd__dlxbp_1 s912 (.D(net406),
    .GATE(clknet_4_6_0_clk),
    .Q(net783),
    .Q_N(net782));
 sky130_fd_sc_hd__dlxtn_2 s913 (.D(net407),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net784));
 sky130_fd_sc_hd__dlxtn_1 s914 (.D(net444),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net785));
 sky130_fd_sc_hd__dlxtn_4 s915 (.D(net445),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net786));
 sky130_fd_sc_hd__dlxtp_1 s916 (.D(net449),
    .GATE(clknet_4_8_0_clk),
    .Q(net787));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s917 (.D(net451),
    .SLEEP_B(clknet_4_10_0_clk),
    .Q(net788));
 sky130_fd_sc_hd__dfxbp_1 s918 (.CLK(clknet_4_9_0_clk),
    .D(net455),
    .Q(net790),
    .Q_N(net789));
 sky130_fd_sc_hd__dfxbp_1 s919 (.CLK(clknet_4_11_0_clk),
    .D(net469),
    .Q(net792),
    .Q_N(net791));
 sky130_fd_sc_hd__dfxtp_4 s920 (.CLK(clknet_4_9_0_clk),
    .D(net472),
    .Q(net793));
 sky130_fd_sc_hd__dfxtp_1 s921 (.CLK(clknet_4_11_0_clk),
    .D(net473),
    .Q(net794));
 sky130_fd_sc_hd__dfxtp_1 s922 (.CLK(clknet_4_9_0_clk),
    .D(net475),
    .Q(net795));
 sky130_fd_sc_hd__dlclkp_1 s923 (.CLK(clknet_4_11_0_clk),
    .GATE(net478),
    .GCLK(net796));
 sky130_fd_sc_hd__dlclkp_2 s924 (.CLK(clknet_4_12_0_clk),
    .GATE(net494),
    .GCLK(net797));
 sky130_fd_sc_hd__dlclkp_4 s925 (.CLK(clknet_4_13_0_clk),
    .GATE(net506),
    .GCLK(net798));
 sky130_fd_sc_hd__dlxbn_1 s926 (.D(net516),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net800),
    .Q_N(net799));
 sky130_fd_sc_hd__dlxbn_2 s927 (.D(net555),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net802),
    .Q_N(net801));
 sky130_fd_sc_hd__dlxbp_1 s928 (.D(net556),
    .GATE(clknet_4_10_0_clk),
    .Q(net804),
    .Q_N(net803));
 sky130_fd_sc_hd__dlxtn_1 s929 (.D(net558),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net805));
 sky130_fd_sc_hd__dlxtn_4 s930 (.D(net559),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net806));
 sky130_fd_sc_hd__dlxtn_1 s931 (.D(net561),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net807));
 sky130_fd_sc_hd__dlxtp_1 s932 (.D(net562),
    .GATE(clknet_4_10_0_clk),
    .Q(net808));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s933 (.D(net563),
    .SLEEP_B(clknet_4_11_0_clk),
    .Q(net809));
 sky130_fd_sc_hd__dfxbp_1 s934 (.CLK(clknet_4_14_0_clk),
    .D(net570),
    .Q(net811),
    .Q_N(net810));
 sky130_fd_sc_hd__dfxbp_1 s935 (.CLK(clknet_4_11_0_clk),
    .D(net573),
    .Q(net813),
    .Q_N(net812));
 sky130_fd_sc_hd__dfxtp_1 s936 (.CLK(clknet_4_11_0_clk),
    .D(net575),
    .Q(net814));
 sky130_fd_sc_hd__dfxtp_1 s937 (.CLK(clknet_4_11_0_clk),
    .D(net576),
    .Q(net815));
 sky130_fd_sc_hd__dfxtp_1 s938 (.CLK(clknet_4_14_0_clk),
    .D(net589),
    .Q(net816));
 sky130_fd_sc_hd__dlclkp_1 s939 (.CLK(clknet_4_14_0_clk),
    .GATE(net594),
    .GCLK(net817));
 sky130_fd_sc_hd__dlclkp_2 s940 (.CLK(clknet_4_14_0_clk),
    .GATE(net603),
    .GCLK(net818));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(in0),
    .X(net165));
 sky130_fd_sc_hd__buf_1 input2 (.A(in1),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(in10),
    .X(net703));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(in11),
    .X(net819));
 sky130_fd_sc_hd__buf_1 input5 (.A(in12),
    .X(net820));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(in13),
    .X(net821));
 sky130_fd_sc_hd__buf_1 input7 (.A(in14),
    .X(net822));
 sky130_fd_sc_hd__buf_2 input8 (.A(in15),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(in16),
    .X(net824));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(in17),
    .X(net825));
 sky130_fd_sc_hd__buf_2 input11 (.A(in18),
    .X(net826));
 sky130_fd_sc_hd__buf_4 input12 (.A(in19),
    .X(net827));
 sky130_fd_sc_hd__buf_4 input13 (.A(in2),
    .X(net828));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(in20),
    .X(net829));
 sky130_fd_sc_hd__buf_4 input15 (.A(in21),
    .X(net830));
 sky130_fd_sc_hd__buf_4 input16 (.A(in22),
    .X(net831));
 sky130_fd_sc_hd__buf_2 input17 (.A(in23),
    .X(net832));
 sky130_fd_sc_hd__buf_2 input18 (.A(in24),
    .X(net833));
 sky130_fd_sc_hd__clkbuf_8 input19 (.A(in25),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(in26),
    .X(net835));
 sky130_fd_sc_hd__buf_2 input21 (.A(in27),
    .X(net836));
 sky130_fd_sc_hd__buf_4 input22 (.A(in28),
    .X(net837));
 sky130_fd_sc_hd__buf_2 input23 (.A(in29),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(in3),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(in30),
    .X(net840));
 sky130_fd_sc_hd__clkbuf_4 input26 (.A(in31),
    .X(net841));
 sky130_fd_sc_hd__buf_4 input27 (.A(in32),
    .X(net842));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(in33),
    .X(net843));
 sky130_fd_sc_hd__clkbuf_8 input29 (.A(in34),
    .X(net844));
 sky130_fd_sc_hd__clkbuf_4 input30 (.A(in35),
    .X(net845));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(in36),
    .X(net846));
 sky130_fd_sc_hd__buf_2 input32 (.A(in37),
    .X(net847));
 sky130_fd_sc_hd__buf_2 input33 (.A(in38),
    .X(net848));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(in39),
    .X(net849));
 sky130_fd_sc_hd__buf_2 input35 (.A(in4),
    .X(net850));
 sky130_fd_sc_hd__dlymetal6s2s_1 input36 (.A(in40),
    .X(net851));
 sky130_fd_sc_hd__clkbuf_4 input37 (.A(in41),
    .X(net852));
 sky130_fd_sc_hd__buf_2 input38 (.A(in42),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_4 input39 (.A(in43),
    .X(net854));
 sky130_fd_sc_hd__buf_1 input40 (.A(in44),
    .X(net855));
 sky130_fd_sc_hd__buf_4 input41 (.A(in45),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(in46),
    .X(net857));
 sky130_fd_sc_hd__clkbuf_4 input43 (.A(in47),
    .X(net858));
 sky130_fd_sc_hd__buf_6 input44 (.A(in48),
    .X(net859));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(in49),
    .X(net860));
 sky130_fd_sc_hd__clkbuf_4 input46 (.A(in5),
    .X(net861));
 sky130_fd_sc_hd__buf_8 input47 (.A(in50),
    .X(net862));
 sky130_fd_sc_hd__clkbuf_4 input48 (.A(in51),
    .X(net863));
 sky130_fd_sc_hd__buf_6 input49 (.A(in52),
    .X(net864));
 sky130_fd_sc_hd__buf_4 input50 (.A(in53),
    .X(net865));
 sky130_fd_sc_hd__buf_2 input51 (.A(in54),
    .X(net866));
 sky130_fd_sc_hd__buf_6 input52 (.A(in55),
    .X(net867));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(in56),
    .X(net868));
 sky130_fd_sc_hd__buf_6 input54 (.A(in57),
    .X(net869));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(in58),
    .X(net870));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(in59),
    .X(net871));
 sky130_fd_sc_hd__clkbuf_4 input57 (.A(in6),
    .X(net872));
 sky130_fd_sc_hd__buf_2 input58 (.A(in60),
    .X(net873));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(in61),
    .X(net874));
 sky130_fd_sc_hd__buf_2 input60 (.A(in7),
    .X(net875));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(in8),
    .X(net876));
 sky130_fd_sc_hd__buf_4 input62 (.A(in9),
    .X(net877));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net878),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(clknet_1_1__leaf_net879),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output65 (.A(net880),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output66 (.A(net960),
    .X(out14));
 sky130_fd_sc_hd__clkbuf_4 output67 (.A(net882),
    .X(out15));
 sky130_fd_sc_hd__clkbuf_4 output68 (.A(net883),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output69 (.A(net884),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output70 (.A(net885),
    .X(out18));
 sky130_fd_sc_hd__clkbuf_4 output71 (.A(net886),
    .X(out19));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net887),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output73 (.A(net888),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output74 (.A(net889),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output75 (.A(net890),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output76 (.A(net891),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output77 (.A(net942),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output78 (.A(net893),
    .X(out25));
 sky130_fd_sc_hd__buf_2 output79 (.A(net894),
    .X(out26));
 sky130_fd_sc_hd__clkbuf_4 output80 (.A(net895),
    .X(out27));
 sky130_fd_sc_hd__clkbuf_4 output81 (.A(net896),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output82 (.A(net897),
    .X(out29));
 sky130_fd_sc_hd__buf_2 output83 (.A(net898),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output84 (.A(net899),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output85 (.A(net946),
    .X(out31));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(clknet_1_1__leaf_net901),
    .X(out32));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(clknet_1_0__leaf_net902),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output88 (.A(net982),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output89 (.A(net904),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(clknet_1_0__leaf_net905),
    .X(out37));
 sky130_fd_sc_hd__clkbuf_4 output91 (.A(net906),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_4 output92 (.A(net907),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output93 (.A(net908),
    .X(out41));
 sky130_fd_sc_hd__clkbuf_4 output94 (.A(net909),
    .X(out42));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(clknet_1_0__leaf_net910),
    .X(out43));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(clknet_1_1__leaf_net911),
    .X(out44));
 sky130_fd_sc_hd__buf_2 output97 (.A(net912),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output98 (.A(net913),
    .X(out46));
 sky130_fd_sc_hd__buf_2 output99 (.A(net952),
    .X(out48));
 sky130_fd_sc_hd__clkbuf_4 output100 (.A(net915),
    .X(out5));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(net916),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output102 (.A(net917),
    .X(out51));
 sky130_fd_sc_hd__buf_2 output103 (.A(net918),
    .X(out52));
 sky130_fd_sc_hd__buf_2 output104 (.A(net919),
    .X(out53));
 sky130_fd_sc_hd__buf_2 output105 (.A(net920),
    .X(out54));
 sky130_fd_sc_hd__buf_2 output106 (.A(net921),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output107 (.A(net990),
    .X(out56));
 sky130_fd_sc_hd__buf_2 output108 (.A(net923),
    .X(out57));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(clknet_1_0__leaf_net924),
    .X(out58));
 sky130_fd_sc_hd__buf_2 output110 (.A(net925),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output111 (.A(net926),
    .X(out60));
 sky130_fd_sc_hd__buf_2 output112 (.A(net927),
    .X(out61));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(net928),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_4 output114 (.A(net929),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output115 (.A(net930),
    .X(out9));
 sky130_fd_sc_hd__buf_4 fanout116 (.A(net909),
    .X(net931));
 sky130_fd_sc_hd__buf_4 fanout117 (.A(net450),
    .X(net932));
 sky130_fd_sc_hd__clkbuf_4 fanout118 (.A(net906),
    .X(net933));
 sky130_fd_sc_hd__clkbuf_4 fanout119 (.A(net441),
    .X(net934));
 sky130_fd_sc_hd__buf_4 fanout120 (.A(net122),
    .X(net935));
 sky130_fd_sc_hd__buf_4 fanout121 (.A(net105),
    .X(net936));
 sky130_fd_sc_hd__buf_2 fanout122 (.A(net340),
    .X(net937));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout123 (.A(net340),
    .X(net938));
 sky130_fd_sc_hd__buf_4 fanout124 (.A(net319),
    .X(net939));
 sky130_fd_sc_hd__clkbuf_2 fanout125 (.A(net319),
    .X(net940));
 sky130_fd_sc_hd__clkbuf_4 fanout126 (.A(net942),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_4 fanout127 (.A(net892),
    .X(net942));
 sky130_fd_sc_hd__clkbuf_4 fanout128 (.A(net919),
    .X(net943));
 sky130_fd_sc_hd__buf_4 fanout129 (.A(net212),
    .X(net944));
 sky130_fd_sc_hd__clkbuf_4 fanout130 (.A(net946),
    .X(net945));
 sky130_fd_sc_hd__clkbuf_4 fanout131 (.A(net947),
    .X(net946));
 sky130_fd_sc_hd__clkbuf_4 fanout132 (.A(net900),
    .X(net947));
 sky130_fd_sc_hd__clkbuf_4 fanout133 (.A(net210),
    .X(net948));
 sky130_fd_sc_hd__buf_4 fanout134 (.A(net101),
    .X(net949));
 sky130_fd_sc_hd__clkbuf_4 fanout135 (.A(net220),
    .X(net950));
 sky130_fd_sc_hd__buf_8 fanout136 (.A(net22),
    .X(net951));
 sky130_fd_sc_hd__clkbuf_4 fanout137 (.A(net914),
    .X(net952));
 sky130_fd_sc_hd__buf_2 fanout138 (.A(net914),
    .X(net953));
 sky130_fd_sc_hd__clkbuf_4 fanout139 (.A(net894),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_4 fanout140 (.A(net956),
    .X(net955));
 sky130_fd_sc_hd__buf_2 fanout141 (.A(net278),
    .X(net956));
 sky130_fd_sc_hd__clkbuf_4 fanout142 (.A(net958),
    .X(net957));
 sky130_fd_sc_hd__buf_2 fanout143 (.A(net959),
    .X(net958));
 sky130_fd_sc_hd__buf_2 fanout144 (.A(net137),
    .X(net959));
 sky130_fd_sc_hd__clkbuf_8 fanout145 (.A(net881),
    .X(net960));
 sky130_fd_sc_hd__buf_4 fanout146 (.A(net88),
    .X(net961));
 sky130_fd_sc_hd__buf_4 fanout147 (.A(net211),
    .X(net962));
 sky130_fd_sc_hd__clkbuf_4 fanout148 (.A(net965),
    .X(net963));
 sky130_fd_sc_hd__clkbuf_4 fanout149 (.A(net965),
    .X(net964));
 sky130_fd_sc_hd__clkbuf_4 fanout150 (.A(net966),
    .X(net965));
 sky130_fd_sc_hd__clkbuf_4 fanout151 (.A(net203),
    .X(net966));
 sky130_fd_sc_hd__buf_4 fanout152 (.A(net199),
    .X(net967));
 sky130_fd_sc_hd__buf_4 fanout153 (.A(net317),
    .X(net968));
 sky130_fd_sc_hd__buf_4 fanout154 (.A(net82),
    .X(net969));
 sky130_fd_sc_hd__buf_8 fanout155 (.A(net971),
    .X(net970));
 sky130_fd_sc_hd__buf_12 fanout156 (.A(net973),
    .X(net971));
 sky130_fd_sc_hd__clkbuf_4 fanout157 (.A(net973),
    .X(net972));
 sky130_fd_sc_hd__buf_6 fanout158 (.A(net17),
    .X(net973));
 sky130_fd_sc_hd__buf_4 fanout159 (.A(net195),
    .X(net974));
 sky130_fd_sc_hd__clkbuf_2 fanout160 (.A(net195),
    .X(net975));
 sky130_fd_sc_hd__buf_2 fanout161 (.A(net977),
    .X(net976));
 sky130_fd_sc_hd__buf_2 fanout162 (.A(net978),
    .X(net977));
 sky130_fd_sc_hd__buf_4 fanout163 (.A(net979),
    .X(net978));
 sky130_fd_sc_hd__buf_4 fanout164 (.A(net189),
    .X(net979));
 sky130_fd_sc_hd__clkbuf_4 fanout165 (.A(net77),
    .X(net980));
 sky130_fd_sc_hd__buf_4 fanout166 (.A(net982),
    .X(net981));
 sky130_fd_sc_hd__buf_4 fanout167 (.A(net903),
    .X(net982));
 sky130_fd_sc_hd__buf_4 fanout168 (.A(net73),
    .X(net983));
 sky130_fd_sc_hd__buf_4 fanout169 (.A(net72),
    .X(net984));
 sky130_fd_sc_hd__clkbuf_4 fanout170 (.A(net794),
    .X(net985));
 sky130_fd_sc_hd__clkbuf_4 fanout171 (.A(net787),
    .X(net986));
 sky130_fd_sc_hd__clkbuf_2 max_cap172 (.A(net768),
    .X(net987));
 sky130_fd_sc_hd__buf_4 fanout173 (.A(net697),
    .X(net988));
 sky130_fd_sc_hd__buf_4 fanout174 (.A(net695),
    .X(net989));
 sky130_fd_sc_hd__buf_12 fanout175 (.A(net922),
    .X(net990));
 sky130_fd_sc_hd__clkbuf_4 fanout176 (.A(net70),
    .X(net991));
 sky130_fd_sc_hd__buf_2 fanout177 (.A(net70),
    .X(net992));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(net69),
    .X(net993));
 sky130_fd_sc_hd__buf_4 fanout179 (.A(net824),
    .X(net994));
 sky130_fd_sc_hd__clkbuf_4 fanout180 (.A(net823),
    .X(net995));
 sky130_fd_sc_hd__clkbuf_4 fanout181 (.A(net822),
    .X(net996));
 sky130_fd_sc_hd__clkbuf_8 fanout182 (.A(net877),
    .X(net997));
 sky130_fd_sc_hd__buf_4 fanout183 (.A(net1001),
    .X(net998));
 sky130_fd_sc_hd__buf_2 fanout184 (.A(net1001),
    .X(net999));
 sky130_fd_sc_hd__buf_4 fanout185 (.A(net1001),
    .X(net1000));
 sky130_fd_sc_hd__clkbuf_4 fanout186 (.A(net876),
    .X(net1001));
 sky130_fd_sc_hd__buf_4 fanout187 (.A(net875),
    .X(net1002));
 sky130_fd_sc_hd__buf_4 fanout188 (.A(net821),
    .X(net1003));
 sky130_fd_sc_hd__buf_4 fanout189 (.A(net872),
    .X(net1004));
 sky130_fd_sc_hd__buf_4 fanout190 (.A(net820),
    .X(net1005));
 sky130_fd_sc_hd__clkbuf_8 fanout191 (.A(net861),
    .X(net1006));
 sky130_fd_sc_hd__clkbuf_4 fanout192 (.A(net855),
    .X(net1007));
 sky130_fd_sc_hd__buf_2 fanout193 (.A(net855),
    .X(net1008));
 sky130_fd_sc_hd__buf_4 fanout194 (.A(net819),
    .X(net1009));
 sky130_fd_sc_hd__clkbuf_4 fanout195 (.A(net851),
    .X(net1010));
 sky130_fd_sc_hd__clkbuf_2 fanout196 (.A(net851),
    .X(net1011));
 sky130_fd_sc_hd__buf_8 fanout197 (.A(net850),
    .X(net1012));
 sky130_fd_sc_hd__clkbuf_8 fanout198 (.A(net848),
    .X(net1013));
 sky130_fd_sc_hd__buf_4 fanout199 (.A(net839),
    .X(net1014));
 sky130_fd_sc_hd__buf_4 fanout200 (.A(net835),
    .X(net1015));
 sky130_fd_sc_hd__buf_4 fanout201 (.A(net176),
    .X(net1016));
 sky130_fd_sc_hd__buf_2 fanout202 (.A(net176),
    .X(net1017));
 sky130_fd_sc_hd__buf_4 fanout203 (.A(net830),
    .X(net1018));
 sky130_fd_sc_hd__buf_4 fanout204 (.A(net829),
    .X(net1019));
 sky130_fd_sc_hd__clkbuf_2 fanout205 (.A(net829),
    .X(net1020));
 sky130_fd_sc_hd__buf_4 fanout206 (.A(net828),
    .X(net1021));
 sky130_fd_sc_hd__buf_4 fanout207 (.A(net1023),
    .X(net1022));
 sky130_fd_sc_hd__clkbuf_8 fanout208 (.A(net826),
    .X(net1023));
 sky130_fd_sc_hd__buf_4 fanout209 (.A(net825),
    .X(net1024));
 sky130_fd_sc_hd__buf_4 fanout210 (.A(net165),
    .X(net1025));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net818 (.A(net818),
    .X(clknet_0_net818));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net818 (.A(clknet_0_net818),
    .X(clknet_1_0__leaf_net818));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net818 (.A(clknet_0_net818),
    .X(clknet_1_1__leaf_net818));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net615 (.A(net615),
    .X(clknet_0_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net615 (.A(clknet_0_net615),
    .X(clknet_1_0__leaf_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net615 (.A(clknet_0_net615),
    .X(clknet_1_1__leaf_net615));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net817 (.A(net817),
    .X(clknet_0_net817));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net817 (.A(clknet_0_net817),
    .X(clknet_1_0__leaf_net817));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net817 (.A(clknet_0_net817),
    .X(clknet_1_1__leaf_net817));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net608 (.A(net608),
    .X(clknet_0_net608));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net608 (.A(clknet_0_net608),
    .X(clknet_1_0__leaf_net608));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net608 (.A(clknet_0_net608),
    .X(clknet_1_1__leaf_net608));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net600 (.A(net600),
    .X(clknet_0_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net600 (.A(clknet_0_net600),
    .X(clknet_1_0__leaf_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net600 (.A(clknet_0_net600),
    .X(clknet_1_1__leaf_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net711 (.A(net711),
    .X(clknet_0_net711));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net711 (.A(clknet_0_net711),
    .X(clknet_1_0__leaf_net711));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net711 (.A(clknet_0_net711),
    .X(clknet_1_1__leaf_net711));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net611 (.A(net611),
    .X(clknet_0_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net611 (.A(clknet_0_net611),
    .X(clknet_1_0__leaf_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net611 (.A(clknet_0_net611),
    .X(clknet_1_1__leaf_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net577 (.A(net577),
    .X(clknet_0_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net577 (.A(clknet_0_net577),
    .X(clknet_1_0__leaf_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net577 (.A(clknet_0_net577),
    .X(clknet_1_1__leaf_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net798 (.A(net798),
    .X(clknet_0_net798));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net798 (.A(clknet_0_net798),
    .X(clknet_1_0__leaf_net798));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net798 (.A(clknet_0_net798),
    .X(clknet_1_1__leaf_net798));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net511 (.A(net511),
    .X(clknet_0_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net511 (.A(clknet_0_net511),
    .X(clknet_1_0__leaf_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net511 (.A(clknet_0_net511),
    .X(clknet_1_1__leaf_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net797 (.A(net797),
    .X(clknet_0_net797));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net797 (.A(clknet_0_net797),
    .X(clknet_1_0__leaf_net797));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net797 (.A(clknet_0_net797),
    .X(clknet_1_1__leaf_net797));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net602 (.A(net602),
    .X(clknet_0_net602));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net602 (.A(clknet_0_net602),
    .X(clknet_1_0__leaf_net602));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net602 (.A(clknet_0_net602),
    .X(clknet_1_1__leaf_net602));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net495 (.A(net495),
    .X(clknet_0_net495));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net495 (.A(clknet_0_net495),
    .X(clknet_1_0__leaf_net495));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net495 (.A(clknet_0_net495),
    .X(clknet_1_1__leaf_net495));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net502 (.A(net502),
    .X(clknet_0_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net502 (.A(clknet_0_net502),
    .X(clknet_1_0__leaf_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net502 (.A(clknet_0_net502),
    .X(clknet_1_1__leaf_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net796 (.A(net796),
    .X(clknet_0_net796));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net796 (.A(clknet_0_net796),
    .X(clknet_1_0__leaf_net796));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net796 (.A(clknet_0_net796),
    .X(clknet_1_1__leaf_net796));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net777 (.A(net777),
    .X(clknet_0_net777));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net777 (.A(clknet_0_net777),
    .X(clknet_1_0__leaf_net777));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net777 (.A(clknet_0_net777),
    .X(clknet_1_1__leaf_net777));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net398 (.A(net398),
    .X(clknet_0_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_0__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_1__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net610 (.A(net610),
    .X(clknet_0_net610));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net610 (.A(clknet_0_net610),
    .X(clknet_1_0__leaf_net610));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net610 (.A(clknet_0_net610),
    .X(clknet_1_1__leaf_net610));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net420 (.A(net420),
    .X(clknet_0_net420));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net420 (.A(clknet_0_net420),
    .X(clknet_1_0__leaf_net420));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net420 (.A(clknet_0_net420),
    .X(clknet_1_1__leaf_net420));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net391 (.A(net391),
    .X(clknet_0_net391));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net391 (.A(clknet_0_net391),
    .X(clknet_1_0__leaf_net391));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net391 (.A(clknet_0_net391),
    .X(clknet_1_1__leaf_net391));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net389 (.A(net389),
    .X(clknet_0_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_0__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_1__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net776 (.A(net776),
    .X(clknet_0_net776));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net776 (.A(clknet_0_net776),
    .X(clknet_1_0__leaf_net776));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net776 (.A(clknet_0_net776),
    .X(clknet_1_1__leaf_net776));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net775 (.A(net775),
    .X(clknet_0_net775));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net775 (.A(clknet_0_net775),
    .X(clknet_1_0__leaf_net775));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net775 (.A(clknet_0_net775),
    .X(clknet_1_1__leaf_net775));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net595 (.A(net595),
    .X(clknet_0_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_0__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_1__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net901 (.A(net901),
    .X(clknet_0_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net901 (.A(clknet_0_net901),
    .X(clknet_1_0__leaf_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net901 (.A(clknet_0_net901),
    .X(clknet_1_1__leaf_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net186 (.A(net186),
    .X(clknet_0_net186));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net186 (.A(clknet_0_net186),
    .X(clknet_1_0__leaf_net186));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net186 (.A(clknet_0_net186),
    .X(clknet_1_1__leaf_net186));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net910 (.A(net910),
    .X(clknet_0_net910));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net910 (.A(clknet_0_net910),
    .X(clknet_1_0__leaf_net910));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net910 (.A(clknet_0_net910),
    .X(clknet_1_1__leaf_net910));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net179 (.A(net179),
    .X(clknet_0_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_0__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_1__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net180 (.A(net180),
    .X(clknet_0_net180));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net180 (.A(clknet_0_net180),
    .X(clknet_1_0__leaf_net180));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net180 (.A(clknet_0_net180),
    .X(clknet_1_1__leaf_net180));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net759 (.A(net759),
    .X(clknet_0_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net759 (.A(clknet_0_net759),
    .X(clknet_1_0__leaf_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net759 (.A(clknet_0_net759),
    .X(clknet_1_1__leaf_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net924 (.A(net924),
    .X(clknet_0_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net924 (.A(clknet_0_net924),
    .X(clknet_1_0__leaf_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net924 (.A(clknet_0_net924),
    .X(clknet_1_1__leaf_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net905 (.A(net905),
    .X(clknet_0_net905));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net905 (.A(clknet_0_net905),
    .X(clknet_1_0__leaf_net905));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net905 (.A(clknet_0_net905),
    .X(clknet_1_1__leaf_net905));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net177 (.A(net177),
    .X(clknet_0_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net177 (.A(clknet_0_net177),
    .X(clknet_1_0__leaf_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net177 (.A(clknet_0_net177),
    .X(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net902 (.A(net902),
    .X(clknet_0_net902));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net902 (.A(clknet_0_net902),
    .X(clknet_1_0__leaf_net902));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net902 (.A(clknet_0_net902),
    .X(clknet_1_1__leaf_net902));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net709 (.A(net709),
    .X(clknet_0_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net709 (.A(clknet_0_net709),
    .X(clknet_1_0__leaf_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net709 (.A(clknet_0_net709),
    .X(clknet_1_1__leaf_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net758 (.A(net758),
    .X(clknet_0_net758));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net758 (.A(clknet_0_net758),
    .X(clknet_1_0__leaf_net758));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net758 (.A(clknet_0_net758),
    .X(clknet_1_1__leaf_net758));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net281 (.A(net281),
    .X(clknet_0_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net281 (.A(clknet_0_net281),
    .X(clknet_1_0__leaf_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net281 (.A(clknet_0_net281),
    .X(clknet_1_1__leaf_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net911 (.A(net911),
    .X(clknet_0_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net911 (.A(clknet_0_net911),
    .X(clknet_1_0__leaf_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net911 (.A(clknet_0_net911),
    .X(clknet_1_1__leaf_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net276 (.A(net276),
    .X(clknet_0_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net276 (.A(clknet_0_net276),
    .X(clknet_1_0__leaf_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net276 (.A(clknet_0_net276),
    .X(clknet_1_1__leaf_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net170 (.A(net170),
    .X(clknet_0_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net170 (.A(clknet_0_net170),
    .X(clknet_1_0__leaf_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net170 (.A(clknet_0_net170),
    .X(clknet_1_1__leaf_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net744 (.A(net744),
    .X(clknet_0_net744));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net744 (.A(clknet_0_net744),
    .X(clknet_1_0__leaf_net744));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net744 (.A(clknet_0_net744),
    .X(clknet_1_1__leaf_net744));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net532 (.A(net532),
    .X(clknet_0_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net532 (.A(clknet_0_net532),
    .X(clknet_1_0__leaf_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net532 (.A(clknet_0_net532),
    .X(clknet_1_1__leaf_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net879 (.A(net879),
    .X(clknet_0_net879));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net879 (.A(clknet_0_net879),
    .X(clknet_1_0__leaf_net879));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net879 (.A(clknet_0_net879),
    .X(clknet_1_1__leaf_net879));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net710 (.A(net710),
    .X(clknet_0_net710));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net710 (.A(clknet_0_net710),
    .X(clknet_1_0__leaf_net710));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net710 (.A(clknet_0_net710),
    .X(clknet_1_1__leaf_net710));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net19),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net1026),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net19),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net24),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net21),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net155),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net1031),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net1031),
    .X(net1033));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer9 (.A(net41),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net1078),
    .X(net1035));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer11 (.A(net1035),
    .X(net1036));
 sky130_fd_sc_hd__a41o_1 clone12 (.A1(net28),
    .A2(net871),
    .A3(net42),
    .A4(net856),
    .B1(net1073),
    .X(net1037));
 sky130_fd_sc_hd__clkbuf_1 clone13 (.A(net1077),
    .X(net1038));
 sky130_fd_sc_hd__clkbuf_1 clone14 (.A(net22),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net22),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net154),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net23),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net1042),
    .X(net1043));
 sky130_fd_sc_hd__clkbuf_1 clone19 (.A(net973),
    .X(net1044));
 sky130_fd_sc_hd__clkbuf_1 clone20 (.A(net971),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net799),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net816),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net757),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net753),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net727),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net792),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net346),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net453),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net699),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net921),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net764),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net772),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net805),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net735),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net435),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net663),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net432),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net800),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net809),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net769),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net747),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net770),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net986),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net734),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net704),
    .X(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A2 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_A1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A0 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_B (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_X (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_S0 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_B1_N (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_B1_N (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_X (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A2 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A1 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A4 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A2 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A2 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_S0 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_B (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_Y (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A4 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A0 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A3 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A3 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_X (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A3 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A3 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_X (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A3 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A3 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_X (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A0 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A4 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A0 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A3 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_X (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A3 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_X (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A3 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_X (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A0 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_SCD (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_B1_N (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B1_N (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_B1_N (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_X (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A0 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A3 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A3 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_X (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_S0 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A0 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S0 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A3 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_X (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A0 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A3 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S0 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_SCD (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A4 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_X (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_S0 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_X (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A3 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A0 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A4 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_X (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S0 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_X (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_X (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A0 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_SCD (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_X (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A0 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S0 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A3 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_X (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A0 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A0 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_X (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A3 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A3 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A3 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_X (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A3 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A4 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_X (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_S0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_D (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_X (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A4 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_X (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A4 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_Q_N (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S0 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_S1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A3 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_X (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A0 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_X (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A3 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A3 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_Q_N (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_X (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S0 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A3 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer16_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_S1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A3 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_X (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_X (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_S1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_Q_N (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A4 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A3 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_X (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A4 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A3 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A3 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_X (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A3 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A4 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B1_N (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A3 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_X (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A4 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_X (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A0 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_X (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_X (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A0 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A3 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_S0 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_S0 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_X (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A3 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_S1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B1_N (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_X (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A0 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A3 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_X (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A0 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_X (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_A2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_X (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_S0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A0 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_X (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A2 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A2 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_B1_N (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_A1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A4 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A0 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_X (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_B1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_X (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A3 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A0 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_X (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A3 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A0 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A3 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B1_N (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_X (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A3 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A0 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A3 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_S0 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S0 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_X (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_X (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S0 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S0 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_X (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A0 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S0 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_X (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A0 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_S0 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A3 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A3 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A3 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_B1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_X (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A0 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A0 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_X (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A0 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A4 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_X (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S0 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A0 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A0 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_S1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A2 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_X (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A0 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_S1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A3 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A2 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_X (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A2 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_S1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A3 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A3 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_X (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A2 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_X (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A3 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B1_N (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A4 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_X (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A3 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_X (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A3 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_X (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A0 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_X (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A0 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_RESET_B (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A0 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_X (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer17_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A2 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_X (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A0 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A3 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A3 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A3 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A3 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_X (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_S0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A4 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_Q_N (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_Q (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A0 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_X (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A0 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_S0 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_X (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A3 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_X (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A3 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A3 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_X (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A0 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A2 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A2 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A3 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A0 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_X (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_B1_N (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_X (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A3 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A3 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A3 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A0 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_X (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A0 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A3 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_X (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A0 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S0 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A0 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S0 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_X (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A3 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A3 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_X (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S0 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A3 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_X (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A0 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S0 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S0 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_X (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S0 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A0 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S0 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_X (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone12_A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_A3 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_X (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_X (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_X (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A0 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_SCD (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_B1_N (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_X (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A3 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A3 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_B (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_X (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_X (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A3 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A3 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A0 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A3 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A3 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_B1_N (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_Y (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A3 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_RESET_B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A3 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_X (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S0 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A0 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_X (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A0 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A3 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_Y (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A0 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_X (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_X (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A0 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_SET_B (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A0 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_S0 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A2 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A2 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A2 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_X (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A0 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A3 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A0 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_X (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A0 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A3 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A2 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A2 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A3 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_S0 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_X (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A2 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_D (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_X (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_X (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A0 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_B1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_X (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A0 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A2 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_X (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A0 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A3 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_X (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A0 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A2 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_X (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A3 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_X (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A3 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_SCE (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A4 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_X (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A2 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A3 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_X (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A0 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_RESET_B (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_SCD (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_RESET_B (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_X (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A2 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A3 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_X (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A3 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A0 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A2 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_S0 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_X (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold27_A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A3 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S0 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S0 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A3 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_Q_N (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A0 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A2 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A2 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_Q (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_X (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A0 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_S0 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A3 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A3 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A0 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A3 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A2 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A3 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_X (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A4 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A1 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer10_A (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_X (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S0 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A0 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A2 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A0 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A0 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_X (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_SCD (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_B1_N (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_X (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_X (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A2 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_X (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A1 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A2 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A3 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_S1 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A4 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_X (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S1 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A3 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A1 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A1 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A1 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_X (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A0 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_SCD (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_S0 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_X (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A3 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_S0 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A3 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_Q_N (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A0 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A3 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_X (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A1 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_S0 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A0 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A3 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A3 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_S0 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_X (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A0 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A3 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_SCE (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A3 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_X (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A0 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_X (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A3 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_X (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A3 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A3 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_SCD (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A3 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A4 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_X (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A0 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_X (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A0 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A2 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S0 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A1 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_RESET_B (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_X (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A0 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S1 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A2 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_X (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A3 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_X (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A0 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A1 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_X (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A0 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_X (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_X (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A0 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_S0 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_B1_N (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_X (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A0 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_X (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A0 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A2 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_X (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A0 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_Q (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A0 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A2 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_B1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_X (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A0 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A0 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A3 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_SCD (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_X (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A2 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A2 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_X (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A1 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A0 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_X (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A2 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A3 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A0 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A3 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A3 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_X (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_D (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_X (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_B1_N (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_Y (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_S0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A3 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A3 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_D (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_X (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_Q (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S0 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S0 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_S0 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_S0 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_S0 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A3 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_Q_N (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_SCE (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_S0 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_X (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_Q_N (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S0 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A3 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S0 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A3 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A3 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A3 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_SET_B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B1_N (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_X (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_Q (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S0 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S0 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A2 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S0 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A3 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A3 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_Q (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_S0 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_Q (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_Q (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S0 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S0 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S0 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A4 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A4 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S0 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_B1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold29_A (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_Q (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S0 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S0 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S0 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_B1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_X (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold45_A (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_Q (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S0 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_S1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_X (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_Q (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A3 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S1 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_S1 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_Q_N (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S1 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S0 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_X (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_S1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_B1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S0 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S0 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge860_Q_N (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A3 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold25_A (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge864_Q (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_S1 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S1 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S1 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_B1 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_Q (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A2 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S0 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_X (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_Q (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S0 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_S1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold34_A (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_Q (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S0 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A3 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_Q (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_S1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S0 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_Q (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S1 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S1 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S0 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_S0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A3 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_S1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_X (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_Q (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S0 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A3 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S0 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_S0 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_B1 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_S1 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_B1 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_B1 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_B1 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_Q (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_S0 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_S0 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A3 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_S0 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge885_Q (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S1 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S0 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_Q (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_S0 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_S0 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold23_A (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_Q (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S1 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S0 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S1 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A3 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_X (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_Q (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S0 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S0 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_Q_N (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_S0 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_Q (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_S0 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap172_A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_Q (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S0 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold32_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_Q (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S0 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_S1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S0 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_Q (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_S1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_S1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_B1_N (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_Y (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_Q (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_S0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A3 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A3 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_S0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A3 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_B1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_S1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_S1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_Q (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_S0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_X (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_Q (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S0 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_S0 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A3 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A3 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_Y (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A3 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_S0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A3 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_X (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_Q (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_S0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_Q (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S0 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_S0 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B1_N (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A3 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_Q_N (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S0 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A3 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_Q (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S0 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A3 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_X (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_SCE (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A3 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B1_N (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_SCE (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_RESET_B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_X (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A2 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_B1_N (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_X (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_SCE (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A3 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_A1 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_A2 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_RESET_B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A3 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A3 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_X (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_X (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A4 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A3 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A4 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_X (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A3 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A3 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_X (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A0 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A3 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A3 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A3 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_A1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A3 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A3 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A1 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A2 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_A (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A2 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A3 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A2 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A3 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_S0 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A3 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A3 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A3 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_A (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A3 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A2 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_B1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_A (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A3 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_S1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A3 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A4 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A4 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_S0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A2 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A3 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A2 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A2 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_B1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A4 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A3 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_A1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A4 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A2 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A0 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A3 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A1 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A2 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A2 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A4 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_S0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A4 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A3 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_A1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A0 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A3 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A4 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_X (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A3 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A2 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A4 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_S0 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A3 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_D (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_B1_N (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A2 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_B1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A4 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A3 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A2 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A3 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A3 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_B1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_A1 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A2 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_B1_N (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A2 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A0 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A2 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A4 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A1 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A2 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B1 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A2 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B1 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_X (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_A2 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_B (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A2 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A0 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A1 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone12_A4 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_B1_N (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_B (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A2 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A3 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A3 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A4 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_A2 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_S1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S0 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A3 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_A2 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A0 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A2 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_X (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_A2 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A2 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A0 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A3 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_S1 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A0 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A0 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A2 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A3 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A2 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A2 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A3 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A3 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A2 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A3 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_B1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A3 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_B1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_X (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_A1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_A2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_B1_N (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_B1_N (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_A2 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A3 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S1 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A0 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_S0 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_X (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A0 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A3 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A1 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A0 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A1 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_A2 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A0 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A2 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A2 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone12_A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_X (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A3 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A0 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A1 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A2 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A4 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_X (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_A1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_RESET_B (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_B1_N (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A1 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A3 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_Q (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A3 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_S0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_A3 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_A1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A3 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A3 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A3 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_B1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_X (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_X (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S0 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_RESET_B (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_X (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A3 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S0 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A3 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A3 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_X (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A2 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_X (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A2 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A3 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_Q (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_S0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A2 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A2 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_SCE (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A2 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A2 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_X (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A2 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_X (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A0 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A2 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A2 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A2 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_X (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_Q (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A3 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_S0 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A2 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_X (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge875_Q (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A3 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_S0 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_Q (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A3 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_S0 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A2 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A2 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_Q (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_Q (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_S0 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_B1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_S0 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_Q (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_X (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A2 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A2 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A2 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_Q (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_X (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_D (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A2 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_X (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S1 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A3 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_Q (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A1 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A2 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_X (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A2 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A2 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_X (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A1 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A3 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_X (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold30_A (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_Q (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_A (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_X (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A3 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A2 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_X (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_Q (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_S1 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S0 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A3 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A2 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A3 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_X (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_X (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_SCE (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A3 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A3 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A3 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_SET_B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A2 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_B1_N (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_X (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_X (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A2 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A0 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A3 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A3 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_RESET_B (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_S0 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_X (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A2 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A3 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_S0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A2 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_X (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S0 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A2 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A2 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_X (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A3 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A4 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_SCE (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A4 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_S0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_X (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A3 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A4 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A4 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_B1_N (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A3 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_X (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A3 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A3 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A3 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_S1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_X (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A0 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A3 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_A1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_SCE (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A3 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A2 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A4 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A0 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A2 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_X (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_S1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A3 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A3 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_X (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_S0 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_SET_B (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A4 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_B1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_S1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_X (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A2 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A2 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_X (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_S0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A3 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A3 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A2 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B1_N (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A3 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_B1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A3 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A2 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_X (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_S1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A3 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S0 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S0 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_SET_B (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A2 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_B1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_X (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_SCE (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A3 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_B1_N (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A3 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A3 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_X (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A0 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_B1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A0 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A2 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_SCD (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_X (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A2 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A2 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A4 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A3 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A2 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S0 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_X (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S0 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A0 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A3 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A2 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A0 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A2 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A3 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A4 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_B1 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_B1_N (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_X (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S0 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A3 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_S1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A3 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_X (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A3 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_B1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_B1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_B1_N (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_S0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_S1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A2 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A4 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_B1_N (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_B1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_X (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S0 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A3 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_X (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A4 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_S0 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_S1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_S0 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A3 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_S1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_SCD (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_B1_N (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_X (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S0 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_S0 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S0 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A3 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_X (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_S0 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A3 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A0 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_X (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_S0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_B1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_X (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_S0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_S0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A3 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A4 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_X (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A4 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_X (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A4 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B1_N (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_S1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_B1_N (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_X (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_S0 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_B1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B1_N (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_B1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_D (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_SCE (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_B1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_B1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A3 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A3 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_X (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_S0 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B1_N (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_B1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_X (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A3 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_S1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A0 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_X (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_S1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S0 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A4 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_B1_N (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A4 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_X (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_S0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A4 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A3 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A3 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A3 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A4 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_X (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A2 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S1 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A1 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A4 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A2 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S0 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A3 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A4 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_RESET_B (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A3 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone20_A (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_X (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_S0 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_S0 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A4 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_A4 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_X (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_S1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A3 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_B1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_B1_N (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A3 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_S0 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A3 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_A1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_X (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_S0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_B1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_B1_N (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A2 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A2 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A2 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_X (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A3 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_S0 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A3 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A0 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A3 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A2 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_X (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A3 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A2 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A3 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A3 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A3 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_A2 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A4 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_S0 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_X (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S0 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A3 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B1_N (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_A (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_X (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A4 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_B1_N (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_B1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A2 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B1_N (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_S0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_B1_N (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_B1_N (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_X (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_SCE (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_S0 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_S1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_S0 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_X (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A3 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A2 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_B1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_X (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_S0 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A0 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_S0 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A2 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_S1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A4 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_X (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_S1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_B1_N (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_S0 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B1_N (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B1_N (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_X (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_S0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold43_A (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_X (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A3 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_S1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_S1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_B1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_B1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_B1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap172_X (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_X (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A3 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A3 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_B1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A3 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_X (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A3 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A4 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_X (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A4 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S0 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A3 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A1 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_X (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_B1_N (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A3 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A3 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A3 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A0 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B1_N (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B1_N (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A3 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_X (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B1_N (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_S1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A2 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A3 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A2 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_S0 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_X (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S0 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_X (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_S0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A3 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A3 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A3 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_B1_N (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_X (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A3 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_B1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A2 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A2 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B1_N (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B1_N (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_X (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A0 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A0 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A4 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_B1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A3 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_X (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A3 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A3 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_A1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A3 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_S0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_S0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A3 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_X (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A3 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_B1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_S0 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B1_N (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_S1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_S0 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B1_N (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_X (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_S1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_B1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_S1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A4 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_X (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A3 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A3 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_B1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_S0 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_SCE (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_B1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_B1_N (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_X (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_X (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S0 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A2 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A3 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A3 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A3 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_X (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S0 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A4 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_X (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_B1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A3 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B1_N (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_B1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_B1_N (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_X (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A2 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A2 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A3 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_S0 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A2 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_X (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A3 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_S0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_S0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_X (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_B1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A3 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A4 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_RESET_B (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_B1_N (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_B1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_B1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B1_N (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_X (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A3 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_S1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A4 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_X (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_SCD (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A2 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_S0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A4 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A2 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_X (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A2 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A4 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A4 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_B1_N (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_X (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_A1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A3 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A2 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_S0 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_X (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A2 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A0 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_S1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_B1_N (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_X (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A1 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A1 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_S0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A1 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A4 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A3 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_S0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A3 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A4 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_B1 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_X (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_S1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B1_N (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_B1_N (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B1_N (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_B1_N (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_X (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A3 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_S1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A3 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A3 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A3 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A4 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_B1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_X (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_S0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B1_N (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A3 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_X (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_X (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A2 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_S0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A4 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_A2 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_B1_N (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_S1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_X (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A4 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_X (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A0 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A2 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_X (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_A2 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_A2 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A2 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A2 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_S0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_B1_N (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_X (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_B1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_B1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A2 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A4 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_B1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A2 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B1_N (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_X (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A3 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_S0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_X (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A0 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A3 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_S0 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A3 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_S0 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A2 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A2 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_X (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A2 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A2 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A4 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_B1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_B (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge847_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge864_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_SLEEP_B (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s922_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_SLEEP_B (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s929_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s921_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s933_SLEEP_B (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s935_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge877_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s926_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_GATE (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_X (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A2 (.DIODE(clknet_1_1__leaf_net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(clknet_1_1__leaf_net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net879_X (.DIODE(clknet_1_1__leaf_net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer3_X (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A2 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A3 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone12_X (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A2 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_SCE (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_S1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S0 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A2 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_X (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A3 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A2 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_B1 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A1 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_S1 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone19_X (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net961));
 sky130_fd_sc_hd__mux4_1 clone1 (.A0(net862),
    .A1(net860),
    .A2(net840),
    .A3(net871),
    .S0(net990),
    .S1(net858),
    .X(net1071));
 sky130_fd_sc_hd__a41o_1 clone2 (.A1(net28),
    .A2(net871),
    .A3(net42),
    .A4(net856),
    .B1(net1073),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net43),
    .X(net1073));
 sky130_fd_sc_hd__a21bo_1 clone15 (.A1(net0),
    .A2(net860),
    .B1_N(net1),
    .X(net1074));
 sky130_fd_sc_hd__a41o_1 clone16 (.A1(net16),
    .A2(net18),
    .A3(net970),
    .A4(net13),
    .B1(net19),
    .X(net1075));
 sky130_fd_sc_hd__clkbuf_1 clone17 (.A(net922),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net922),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net36),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net36),
    .X(net1079));
 sky130_fd_sc_hd__a31o_1 clone22 (.A1(net6),
    .A2(net951),
    .A3(net8),
    .B1(net970),
    .X(net1080));
 sky130_fd_sc_hd__a21bo_1 clone23 (.A1(net4),
    .A2(net25),
    .B1_N(net856),
    .X(net1081));
 sky130_fd_sc_hd__a41o_1 clone24 (.A1(net884),
    .A2(net951),
    .A3(net664),
    .A4(net754),
    .B1(net755),
    .X(net1082));
 sky130_fd_sc_hd__clkbuf_1 clone25 (.A(net973),
    .X(net1083));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
