module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in3,
    in4,
    in5,
    in6,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out3,
    out4,
    out5,
    out6,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in3;
 input in4;
 input in5;
 input in6;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out3;
 output out4;
 output out5;
 output out6;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net918;
 wire clknet_1_0__leaf_net918;
 wire clknet_1_1__leaf_net918;
 wire clknet_0_net917;
 wire clknet_1_0__leaf_net917;
 wire clknet_1_1__leaf_net917;
 wire clknet_0_net916;
 wire clknet_1_0__leaf_net916;
 wire clknet_1_1__leaf_net916;
 wire clknet_0_net731;
 wire clknet_1_0__leaf_net731;
 wire clknet_1_1__leaf_net731;
 wire clknet_0_net712;
 wire clknet_1_0__leaf_net712;
 wire clknet_1_1__leaf_net712;
 wire clknet_0_net720;
 wire clknet_1_0__leaf_net720;
 wire clknet_1_1__leaf_net720;
 wire clknet_0_net834;
 wire clknet_1_0__leaf_net834;
 wire clknet_1_1__leaf_net834;
 wire clknet_0_net709;
 wire clknet_1_0__leaf_net709;
 wire clknet_1_1__leaf_net709;
 wire clknet_0_net897;
 wire clknet_1_0__leaf_net897;
 wire clknet_1_1__leaf_net897;
 wire clknet_0_net967;
 wire clknet_1_0__leaf_net967;
 wire clknet_1_1__leaf_net967;
 wire clknet_0_net896;
 wire clknet_1_0__leaf_net896;
 wire clknet_1_1__leaf_net896;
 wire clknet_0_net895;
 wire clknet_1_0__leaf_net895;
 wire clknet_1_1__leaf_net895;
 wire clknet_0_net563;
 wire clknet_1_0__leaf_net563;
 wire clknet_1_1__leaf_net563;
 wire clknet_0_net795;
 wire clknet_1_0__leaf_net795;
 wire clknet_1_1__leaf_net795;
 wire clknet_0_net562;
 wire clknet_1_0__leaf_net562;
 wire clknet_1_1__leaf_net562;
 wire clknet_0_net876;
 wire clknet_1_0__leaf_net876;
 wire clknet_1_1__leaf_net876;
 wire clknet_0_net473;
 wire clknet_1_0__leaf_net473;
 wire clknet_1_1__leaf_net473;
 wire clknet_0_net597;
 wire clknet_1_0__leaf_net597;
 wire clknet_1_1__leaf_net597;
 wire clknet_0_net471;
 wire clknet_1_0__leaf_net471;
 wire clknet_1_1__leaf_net471;
 wire clknet_0_net593;
 wire clknet_1_0__leaf_net593;
 wire clknet_1_1__leaf_net593;
 wire clknet_0_net875;
 wire clknet_1_0__leaf_net875;
 wire clknet_1_1__leaf_net875;
 wire clknet_0_net966;
 wire clknet_1_0__leaf_net966;
 wire clknet_1_1__leaf_net966;
 wire clknet_0_net721;
 wire clknet_1_0__leaf_net721;
 wire clknet_1_1__leaf_net721;
 wire clknet_0_net833;
 wire clknet_1_0__leaf_net833;
 wire clknet_1_1__leaf_net833;
 wire clknet_0_net874;
 wire clknet_1_0__leaf_net874;
 wire clknet_1_1__leaf_net874;
 wire clknet_0_net622;
 wire clknet_1_0__leaf_net622;
 wire clknet_1_1__leaf_net622;
 wire clknet_0_net856;
 wire clknet_1_0__leaf_net856;
 wire clknet_1_1__leaf_net856;
 wire clknet_0_net352;
 wire clknet_1_0__leaf_net352;
 wire clknet_1_1__leaf_net352;
 wire clknet_0_net346;
 wire clknet_1_0__leaf_net346;
 wire clknet_1_1__leaf_net346;
 wire clknet_0_net855;
 wire clknet_1_0__leaf_net855;
 wire clknet_1_1__leaf_net855;
 wire clknet_0_net854;
 wire clknet_1_0__leaf_net854;
 wire clknet_1_1__leaf_net854;
 wire clknet_0_net227;
 wire clknet_1_0__leaf_net227;
 wire clknet_1_1__leaf_net227;
 wire clknet_0_net958;
 wire clknet_1_0__leaf_net958;
 wire clknet_1_1__leaf_net958;
 wire clknet_0_net229;
 wire clknet_1_0__leaf_net229;
 wire clknet_1_1__leaf_net229;
 wire clknet_0_net228;
 wire clknet_1_0__leaf_net228;
 wire clknet_1_1__leaf_net228;
 wire clknet_0_net222;
 wire clknet_1_0__leaf_net222;
 wire clknet_1_1__leaf_net222;
 wire clknet_0_net798;
 wire clknet_1_0__leaf_net798;
 wire clknet_1_1__leaf_net798;
 wire clknet_0_net215;
 wire clknet_1_0__leaf_net215;
 wire clknet_1_1__leaf_net215;
 wire clknet_0_net91;
 wire clknet_1_0__leaf_net91;
 wire clknet_1_1__leaf_net91;
 wire clknet_0_net97;
 wire clknet_1_0__leaf_net97;
 wire clknet_1_1__leaf_net97;
 wire clknet_0_net96;
 wire clknet_1_0__leaf_net96;
 wire clknet_1_1__leaf_net96;
 wire clknet_0_net232;
 wire clknet_1_0__leaf_net232;
 wire clknet_1_1__leaf_net232;
 wire clknet_0_net95;
 wire clknet_1_0__leaf_net95;
 wire clknet_1_1__leaf_net95;
 wire clknet_0_net94;
 wire clknet_1_0__leaf_net94;
 wire clknet_1_1__leaf_net94;
 wire clknet_0_net98;
 wire clknet_1_0__leaf_net98;
 wire clknet_1_1__leaf_net98;
 wire clknet_0_net102;
 wire clknet_1_0__leaf_net102;
 wire clknet_1_1__leaf_net102;
 wire clknet_0_net797;
 wire clknet_1_0__leaf_net797;
 wire clknet_1_1__leaf_net797;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;

 sky130_fd_sc_hd__and3_2 c100 (.A(net68),
    .B(net52),
    .C(net1001),
    .X(net73));
 sky130_fd_sc_hd__a2111o_1 c101 (.A1(net66),
    .A2(net68),
    .B1(net991),
    .C1(net43),
    .D1(net6),
    .X(net74));
 sky130_fd_sc_hd__a2111o_2 c102 (.A1(net1084),
    .A2(net69),
    .B1(net57),
    .C1(net67),
    .D1(net28),
    .X(net75));
 sky130_fd_sc_hd__and2_0 c103 (.A(net64),
    .B(net1001),
    .X(net76));
 sky130_fd_sc_hd__and3_1 c104 (.A(net55),
    .B(net74),
    .C(net76),
    .X(net77));
 sky130_fd_sc_hd__and3_1 c105 (.A(net75),
    .B(net32),
    .C(net1022),
    .X(net78));
 sky130_fd_sc_hd__and2_1 c106 (.A(net74),
    .B(net941),
    .X(net79));
 sky130_fd_sc_hd__and2_0 c107 (.A(net52),
    .B(net76),
    .X(net80));
 sky130_fd_sc_hd__a2111o_4 c108 (.A1(net43),
    .A2(net74),
    .B1(net1022),
    .C1(net991),
    .D1(net1001),
    .X(net81));
 sky130_fd_sc_hd__and3_1 c109 (.A(net76),
    .B(net80),
    .C(net1001),
    .X(net82));
 sky130_fd_sc_hd__and3_1 c110 (.A(net944),
    .B(net49),
    .C(net20),
    .X(net83));
 sky130_fd_sc_hd__or4bb_4 c111 (.A(net928),
    .B(net20),
    .C_N(net69),
    .D_N(net1002),
    .X(net84));
 sky130_fd_sc_hd__a2111o_4 c112 (.A1(net945),
    .A2(net928),
    .B1(net991),
    .C1(net1062),
    .D1(net83),
    .X(net85));
 sky130_fd_sc_hd__and3_2 c113 (.A(net83),
    .B(net10),
    .C(net1002),
    .X(net86));
 sky130_fd_sc_hd__and3_1 c114 (.A(net72),
    .B(net83),
    .C(net1048),
    .X(net87));
 sky130_fd_sc_hd__and3_1 c115 (.A(net3),
    .B(net20),
    .C(net69),
    .X(net88));
 sky130_fd_sc_hd__a2111o_4 c116 (.A1(net13),
    .A2(net87),
    .B1(net991),
    .C1(net1002),
    .D1(net85),
    .X(net89));
 sky130_fd_sc_hd__and3_1 c117 (.A(net88),
    .B(net85),
    .C(net1002),
    .X(net90));
 sky130_fd_sc_hd__buf_1 c118 (.A(clknet_1_1__leaf_net798),
    .X(net91));
 sky130_fd_sc_hd__and3_2 c119 (.A(net80),
    .B(net86),
    .C(net1022),
    .X(net92));
 sky130_fd_sc_hd__or4bb_1 c120 (.A(net20),
    .B(net77),
    .C_N(net89),
    .D_N(net1158),
    .X(net93));
 sky130_fd_sc_hd__and3_1 c121 (.A(clknet_1_0__leaf_net91),
    .B(net83),
    .C(net86),
    .X(net94));
 sky130_fd_sc_hd__a2111o_1 c122 (.A1(net87),
    .A2(net992),
    .B1(net85),
    .C1(clknet_1_1__leaf_net91),
    .D1(net88),
    .X(net95));
 sky130_fd_sc_hd__a2111o_1 c123 (.A1(clknet_1_0__leaf_net94),
    .A2(net88),
    .B1(net85),
    .C1(clknet_1_0__leaf_net91),
    .D1(net1041),
    .X(net96));
 sky130_fd_sc_hd__and3_1 c124 (.A(net90),
    .B(net50),
    .C(clknet_1_1__leaf_net91),
    .X(net97));
 sky130_fd_sc_hd__a2111o_1 c125 (.A1(net69),
    .A2(clknet_1_1__leaf_net94),
    .B1(net992),
    .C1(net10),
    .D1(net86),
    .X(net98));
 sky130_fd_sc_hd__mux4_1 c126 (.A0(net38),
    .A1(clknet_1_0__leaf_net97),
    .A2(net89),
    .A3(clknet_1_0__leaf_net96),
    .S0(net1037),
    .S1(net84),
    .X(net99));
 sky130_fd_sc_hd__mux4_1 c127 (.A0(clknet_1_0__leaf_net97),
    .A1(clknet_1_1__leaf_net91),
    .A2(net87),
    .A3(net38),
    .S0(clknet_1_1__leaf_net98),
    .S1(net848),
    .X(net100));
 sky130_fd_sc_hd__a2111o_1 c128 (.A1(net90),
    .A2(net85),
    .B1(clknet_1_0__leaf_net95),
    .D1(net847),
    .X(net101));
 sky130_fd_sc_hd__or4bb_1 c129 (.A(clknet_1_0__leaf_net98),
    .B(net13),
    .C_N(net764),
    .D_N(net847),
    .X(net102));
 sky130_fd_sc_hd__a2111o_1 c130 (.A1(net992),
    .A2(net944),
    .B1(net90),
    .C1(clknet_1_0__leaf_net102),
    .D1(net763),
    .X(net103));
 sky130_fd_sc_hd__sdfbbn_1 c131 (.CLK_N(clknet_4_4_0_clk),
    .D(clknet_1_1__leaf_net102),
    .RESET_B(net83),
    .SCD(clknet_1_1__leaf_net97),
    .SCE(net89),
    .SET_B(net849),
    .Q(net105),
    .Q_N(net104));
 sky130_fd_sc_hd__and3_4 c132 (.A(net1047),
    .B(net1051),
    .C(net951),
    .X(net106));
 sky130_fd_sc_hd__and2_4 c133 (.A(net930),
    .B(net1054),
    .X(net107));
 sky130_fd_sc_hd__and2_4 c134 (.A(net1057),
    .B(net1058),
    .X(net959));
 sky130_fd_sc_hd__and2_1 c135 (.A(net1059),
    .B(net949),
    .X(net108));
 sky130_fd_sc_hd__and2_4 c136 (.A(net106),
    .B(net1044),
    .X(net109));
 sky130_fd_sc_hd__and2_4 c137 (.A(net1057),
    .B(net951),
    .X(net110));
 sky130_fd_sc_hd__and2_4 c138 (.A(net1044),
    .B(net939),
    .X(net111));
 sky130_fd_sc_hd__and2_4 c139 (.A(net1042),
    .B(net106),
    .X(net112));
 sky130_fd_sc_hd__and2_2 c140 (.A(net949),
    .B(net1042),
    .X(net113));
 sky130_fd_sc_hd__and2_4 c141 (.A(net109),
    .B(net107),
    .X(net114));
 sky130_fd_sc_hd__and3_4 c142 (.A(net1042),
    .B(net1054),
    .C(net1060),
    .X(net115));
 sky130_fd_sc_hd__and2_4 c143 (.A(net115),
    .B(net1043),
    .X(net116));
 sky130_fd_sc_hd__and2_4 c144 (.A(net116),
    .B(net108),
    .X(net117));
 sky130_fd_sc_hd__and2_4 c145 (.A(net114),
    .B(net116),
    .X(net118));
 sky130_fd_sc_hd__and2_2 c146 (.A(net928),
    .B(net933),
    .X(net119));
 sky130_fd_sc_hd__and2_4 c147 (.A(net111),
    .B(net1042),
    .X(net120));
 sky130_fd_sc_hd__and2_2 c148 (.A(net1126),
    .B(net117),
    .X(net121));
 sky130_fd_sc_hd__and2_2 c149 (.A(net113),
    .B(net1026),
    .X(net122));
 sky130_fd_sc_hd__and2_4 c150 (.A(net109),
    .B(net117),
    .X(net970));
 sky130_fd_sc_hd__mux4_2 c151 (.A0(net118),
    .A1(net117),
    .A2(net1024),
    .A3(net1026),
    .S0(net1042),
    .S1(net119),
    .X(net123));
 sky130_fd_sc_hd__a2111o_4 c152 (.A1(net1060),
    .A2(net123),
    .B1(net1024),
    .C1(net1042),
    .D1(net1044),
    .X(net124));
 sky130_fd_sc_hd__a2111o_4 c153 (.A1(net124),
    .A2(net119),
    .B1(net1024),
    .C1(net970),
    .D1(net1042),
    .X(net125));
 sky130_fd_sc_hd__and2_1 c154 (.A(net114),
    .B(net1038),
    .X(net126));
 sky130_fd_sc_hd__and2_2 c155 (.A(net117),
    .B(net14),
    .X(net127));
 sky130_fd_sc_hd__and2_1 c156 (.A(net106),
    .B(net0),
    .X(net128));
 sky130_fd_sc_hd__and2_1 c157 (.A(net941),
    .B(net1),
    .X(net129));
 sky130_fd_sc_hd__and2_1 c158 (.A(net1059),
    .B(net129),
    .X(net130));
 sky130_fd_sc_hd__and2_1 c159 (.A(net127),
    .B(net119),
    .X(net131));
 sky130_fd_sc_hd__and2_4 c160 (.A(net1051),
    .B(net1038),
    .X(net132));
 sky130_fd_sc_hd__and2_1 c161 (.A(net128),
    .B(net9),
    .X(net133));
 sky130_fd_sc_hd__and2_2 c162 (.A(net1025),
    .B(net126),
    .X(net134));
 sky130_fd_sc_hd__and2_4 c163 (.A(net119),
    .B(net126),
    .X(net135));
 sky130_fd_sc_hd__and2_2 c164 (.A(net129),
    .B(net131),
    .X(net136));
 sky130_fd_sc_hd__and2_1 c165 (.A(net1058),
    .B(net119),
    .X(net137));
 sky130_fd_sc_hd__and3_2 c166 (.A(net941),
    .B(net951),
    .C(net134),
    .X(net138));
 sky130_fd_sc_hd__mux4_2 c167 (.A0(net941),
    .A1(net136),
    .A2(net135),
    .A3(net5),
    .S0(net138),
    .S1(net1018),
    .X(net139));
 sky130_fd_sc_hd__mux4_2 c168 (.A0(net129),
    .A1(net134),
    .A2(net1000),
    .A3(net1018),
    .S0(net1038),
    .S1(net114),
    .X(net140));
 sky130_fd_sc_hd__and3_2 c169 (.A(net136),
    .B(net126),
    .C(net970),
    .X(net141));
 sky130_fd_sc_hd__and2_4 c170 (.A(net130),
    .B(net140),
    .X(net142));
 sky130_fd_sc_hd__a2111o_4 c171 (.A1(net137),
    .A2(net140),
    .B1(net1060),
    .C1(net941),
    .D1(net1126),
    .X(net143));
 sky130_fd_sc_hd__and2_4 c172 (.A(net138),
    .B(net137),
    .X(net144));
 sky130_fd_sc_hd__and2_2 c173 (.A(net1062),
    .B(net137),
    .X(net145));
 sky130_fd_sc_hd__and2_2 c174 (.A(net15),
    .B(net136),
    .X(net146));
 sky130_fd_sc_hd__mux4_2 c175 (.A0(net146),
    .A1(net145),
    .A2(net142),
    .A3(net136),
    .S0(net1018),
    .S1(net1000),
    .X(net147));
 sky130_fd_sc_hd__and3_2 c176 (.A(net1011),
    .B(net111),
    .C(net121),
    .X(net148));
 sky130_fd_sc_hd__or4bb_2 c177 (.A(net1052),
    .B(net109),
    .C_N(net1041),
    .D_N(net28),
    .X(net149));
 sky130_fd_sc_hd__and2_2 c178 (.A(net5),
    .B(net148),
    .X(net150));
 sky130_fd_sc_hd__and2_2 c179 (.A(net35),
    .B(net10),
    .X(net151));
 sky130_fd_sc_hd__and3_2 c180 (.A(net8),
    .B(net106),
    .C(net138),
    .X(net152));
 sky130_fd_sc_hd__and3_2 c181 (.A(net125),
    .B(net149),
    .C(net5),
    .X(net153));
 sky130_fd_sc_hd__a2111o_1 c182 (.A1(net144),
    .A2(net141),
    .B1(net951),
    .C1(net21),
    .D1(net1053),
    .X(net154));
 sky130_fd_sc_hd__and3_2 c183 (.A(net154),
    .B(net151),
    .C(net22),
    .X(net155));
 sky130_fd_sc_hd__or4bb_4 c184 (.A(net151),
    .B(net37),
    .C_N(net1042),
    .D_N(net152),
    .X(net156));
 sky130_fd_sc_hd__a2111o_2 c185 (.A1(net37),
    .A2(net156),
    .B1(net36),
    .C1(net148),
    .D1(net155),
    .X(net157));
 sky130_fd_sc_hd__and3_4 c186 (.A(net928),
    .B(net8),
    .C(net997),
    .X(net158));
 sky130_fd_sc_hd__or4bb_4 c187 (.A(net951),
    .B(net125),
    .C_N(net156),
    .D_N(net152),
    .X(net159));
 sky130_fd_sc_hd__or4bb_4 c188 (.A(net159),
    .B(net150),
    .C_N(net144),
    .D_N(net139),
    .X(net160));
 sky130_fd_sc_hd__a2111o_2 c189 (.A1(net158),
    .A2(net154),
    .B1(net159),
    .C1(net125),
    .D1(net144),
    .X(net161));
 sky130_fd_sc_hd__and2_4 c190 (.A(net5),
    .B(net22),
    .X(net162));
 sky130_fd_sc_hd__or4bb_4 c191 (.A(net156),
    .B(net158),
    .C_N(net134),
    .D_N(net154),
    .X(net163));
 sky130_fd_sc_hd__a2111o_4 c192 (.A1(net160),
    .A2(net131),
    .B1(net109),
    .C1(net163),
    .D1(net1055),
    .X(net164));
 sky130_fd_sc_hd__mux4_2 c193 (.A0(net153),
    .A1(net14),
    .A2(net164),
    .A3(net163),
    .S0(net159),
    .S1(net1018),
    .X(net165));
 sky130_fd_sc_hd__and3_1 c194 (.A(net165),
    .B(net150),
    .C(net163),
    .X(net166));
 sky130_fd_sc_hd__a2111o_2 c195 (.A1(net126),
    .A2(net985),
    .B1(net163),
    .C1(net117),
    .D1(net149),
    .X(net167));
 sky130_fd_sc_hd__a2111o_1 c196 (.A1(net985),
    .A2(net29),
    .B1(net167),
    .C1(net130),
    .D1(net1007),
    .X(net168));
 sky130_fd_sc_hd__a2111o_1 c197 (.A1(net167),
    .A2(net168),
    .B1(net985),
    .C1(net162),
    .D1(net163),
    .X(net169));
 sky130_fd_sc_hd__a2111o_1 c198 (.A1(net135),
    .A2(net37),
    .B1(net46),
    .C1(net985),
    .D1(net157),
    .X(net170));
 sky130_fd_sc_hd__and3_2 c199 (.A(net22),
    .B(net141),
    .C(net124),
    .X(net171));
 sky130_fd_sc_hd__and3_2 c200 (.A(net53),
    .B(net46),
    .C(net50),
    .X(net172));
 sky130_fd_sc_hd__and3_2 c201 (.A(net34),
    .B(net172),
    .C(net111),
    .X(net173));
 sky130_fd_sc_hd__a2111o_4 c202 (.A1(net939),
    .A2(net47),
    .B1(net15),
    .C1(net19),
    .D1(net1025),
    .X(net174));
 sky130_fd_sc_hd__or4bb_4 c203 (.A(net1),
    .B(net1059),
    .C_N(net172),
    .D_N(net1033),
    .X(net175));
 sky130_fd_sc_hd__and3_1 c204 (.A(net170),
    .B(net50),
    .C(net175),
    .X(net176));
 sky130_fd_sc_hd__mux4_1 c205 (.A0(net11),
    .A1(net135),
    .A2(net989),
    .A3(net172),
    .S0(net941),
    .S1(net1051),
    .X(net177));
 sky130_fd_sc_hd__and3_1 c206 (.A(net177),
    .B(net156),
    .C(net175),
    .X(net178));
 sky130_fd_sc_hd__a2111o_1 c207 (.A1(net1054),
    .A2(net53),
    .B1(net57),
    .C1(net60),
    .D1(net170),
    .X(net179));
 sky130_fd_sc_hd__mux4_2 c208 (.A0(net1097),
    .A1(net107),
    .A2(net175),
    .A3(net1018),
    .S0(net171),
    .S1(net1035),
    .X(net180));
 sky130_fd_sc_hd__a2111o_1 c209 (.A1(net59),
    .A2(net138),
    .B1(net149),
    .C1(net985),
    .D1(net996),
    .X(net181));
 sky130_fd_sc_hd__or4bb_1 c210 (.A(net181),
    .B(net177),
    .C_N(net145),
    .D_N(net1041),
    .X(net182));
 sky130_fd_sc_hd__a2111o_1 c211 (.A1(net180),
    .A2(net53),
    .B1(net182),
    .C1(net997),
    .D1(net135),
    .X(net183));
 sky130_fd_sc_hd__a2111o_1 c212 (.A1(net170),
    .A2(net182),
    .B1(net50),
    .C1(net174),
    .D1(net145),
    .X(net184));
 sky130_fd_sc_hd__a2111o_1 c213 (.A1(net14),
    .A2(net184),
    .B1(net172),
    .C1(net171),
    .D1(net985),
    .X(net185));
 sky130_fd_sc_hd__mux4_1 c214 (.A0(net182),
    .A1(net142),
    .A2(net184),
    .A3(net989),
    .S0(net180),
    .S1(net1030),
    .X(net186));
 sky130_fd_sc_hd__a2111o_2 c215 (.A1(net1),
    .A2(net134),
    .B1(net985),
    .C1(net37),
    .D1(net1030),
    .X(net187));
 sky130_fd_sc_hd__mux4_1 c216 (.A0(net184),
    .A1(net170),
    .A2(net138),
    .A3(net59),
    .S0(net15),
    .S1(net983),
    .X(net188));
 sky130_fd_sc_hd__sdfbbn_2 c217 (.CLK_N(clknet_4_1_0_clk),
    .D(net983),
    .RESET_B(net184),
    .SCD(net172),
    .SCE(net1096),
    .SET_B(net1030),
    .Q(net190),
    .Q_N(net189));
 sky130_fd_sc_hd__a2111o_1 c218 (.A1(net149),
    .A2(net181),
    .B1(net983),
    .C1(net989),
    .D1(net1030),
    .X(net191));
 sky130_fd_sc_hd__a2111o_2 c219 (.A1(net145),
    .A2(net983),
    .B1(net54),
    .C1(net189),
    .D1(net1030),
    .X(net192));
 sky130_fd_sc_hd__a2111o_1 c220 (.A1(net46),
    .A2(net989),
    .B1(net172),
    .C1(net189),
    .D1(net1003),
    .X(net193));
 sky130_fd_sc_hd__a2111o_4 c221 (.A1(net941),
    .A2(net176),
    .B1(net73),
    .C1(net1000),
    .D1(net22),
    .X(net194));
 sky130_fd_sc_hd__mux4_1 c222 (.A0(net194),
    .A1(net67),
    .A2(net930),
    .A3(net172),
    .S0(net1000),
    .S1(net1007),
    .X(net195));
 sky130_fd_sc_hd__sdfbbp_1 c223 (.CLK(clknet_4_4_0_clk),
    .D(net82),
    .RESET_B(net71),
    .SCD(net148),
    .SCE(net194),
    .SET_B(net1001),
    .Q(net197),
    .Q_N(net196));
 sky130_fd_sc_hd__a2111o_1 c224 (.A1(net1026),
    .A2(net71),
    .B1(net189),
    .C1(net930),
    .D1(net1035),
    .X(net198));
 sky130_fd_sc_hd__a2111o_1 c225 (.A1(net60),
    .A2(net179),
    .B1(net194),
    .C1(net174),
    .D1(net196),
    .X(net199));
 sky130_fd_sc_hd__mux4_2 c226 (.A0(net193),
    .A1(net164),
    .A2(net1035),
    .A3(net162),
    .S0(net1055),
    .S1(net842),
    .X(net200));
 sky130_fd_sc_hd__mux4_1 c227 (.A0(net930),
    .A1(net194),
    .A2(net1042),
    .A3(net983),
    .S0(net200),
    .S1(net1062),
    .X(net201));
 sky130_fd_sc_hd__a2111o_1 c228 (.A1(net180),
    .A2(net46),
    .B1(net172),
    .C1(net200),
    .D1(net991),
    .X(net202));
 sky130_fd_sc_hd__a2111o_1 c229 (.A1(net179),
    .A2(net194),
    .B1(net200),
    .C1(net991),
    .D1(net180),
    .X(net203));
 sky130_fd_sc_hd__a2111o_1 c230 (.A1(net172),
    .A2(net1083),
    .B1(net158),
    .C1(net2),
    .D1(net134),
    .X(net204));
 sky130_fd_sc_hd__a2111o_1 c231 (.A1(net204),
    .A2(net180),
    .B1(net194),
    .C1(net200),
    .D1(net1147),
    .X(net205));
 sky130_fd_sc_hd__a2111o_1 c232 (.A1(net196),
    .A2(net174),
    .B1(net991),
    .C1(net799),
    .D1(net842),
    .X(net206));
 sky130_fd_sc_hd__a2111o_2 c233 (.A1(net71),
    .A2(net945),
    .B1(net112),
    .C1(net172),
    .D1(net851),
    .X(net207));
 sky130_fd_sc_hd__sdfbbn_1 c234 (.CLK_N(clknet_4_4_0_clk),
    .D(net78),
    .RESET_B(net204),
    .SCD(net200),
    .SCE(net194),
    .SET_B(net799),
    .Q(net209),
    .Q_N(net208));
 sky130_fd_sc_hd__a2111o_2 c235 (.A1(net206),
    .A2(net180),
    .B1(net6),
    .C1(net207),
    .D1(net985),
    .X(net210));
 sky130_fd_sc_hd__mux4_1 c236 (.A0(net194),
    .A1(net989),
    .A2(net174),
    .A3(net1026),
    .S0(net210),
    .S1(net975),
    .X(net211));
 sky130_fd_sc_hd__mux4_2 c237 (.A0(net171),
    .A1(net210),
    .A2(net82),
    .A3(net207),
    .S0(net208),
    .S1(net800),
    .X(net212));
 sky130_fd_sc_hd__a2111o_1 c238 (.A1(net210),
    .A2(net193),
    .B1(net174),
    .C1(net208),
    .D1(net212),
    .X(net213));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net148),
    .A1(net213),
    .A2(net60),
    .A3(net210),
    .S0(net194),
    .S1(net1114),
    .X(net214));
 sky130_fd_sc_hd__mux4_1 c240 (.A0(net202),
    .A1(net60),
    .A2(net180),
    .A3(net77),
    .S0(net210),
    .S1(clknet_1_0__leaf_net798),
    .X(net215));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(net213),
    .A1(net1159),
    .A2(clknet_1_0__leaf_net215),
    .A3(net70),
    .S0(net975),
    .S1(net800),
    .X(net216));
 sky130_fd_sc_hd__mux4_1 c242 (.A0(net124),
    .A1(clknet_1_0__leaf_net215),
    .A2(net75),
    .A3(net1010),
    .S0(net196),
    .S1(net208),
    .X(net217));
 sky130_fd_sc_hd__mux4_1 c243 (.A0(net992),
    .A1(net983),
    .A2(net89),
    .A3(net997),
    .S0(net92),
    .S1(clknet_1_0__leaf_net96),
    .X(net218));
 sky130_fd_sc_hd__mux4_1 c244 (.A0(clknet_1_1__leaf_net215),
    .A1(net152),
    .A2(clknet_1_0__leaf_net96),
    .A3(net983),
    .S0(net1025),
    .S1(net853),
    .X(net219));
 sky130_fd_sc_hd__mux4_1 c245 (.A0(net89),
    .A1(net197),
    .A2(net928),
    .A3(net1002),
    .S0(clknet_1_1__leaf_net798),
    .S1(net853),
    .X(net220));
 sky130_fd_sc_hd__mux4_1 c246 (.A0(net77),
    .A1(net160),
    .A2(net928),
    .A3(net89),
    .S0(net848),
    .S1(net850),
    .X(net221));
 sky130_fd_sc_hd__mux4_1 c247 (.A0(net1097),
    .A1(net50),
    .A2(net118),
    .A3(net57),
    .S0(net853),
    .S1(clknet_1_1__leaf_net854),
    .X(net222));
 sky130_fd_sc_hd__mux4_1 c248 (.A0(net1059),
    .A1(net197),
    .A2(net89),
    .A3(net848),
    .S0(net852),
    .S1(clknet_1_0__leaf_net854),
    .X(net223));
 sky130_fd_sc_hd__mux4_1 c249 (.A0(clknet_1_0__leaf_net95),
    .A1(net209),
    .A2(net89),
    .A3(net1010),
    .S0(net1126),
    .S1(net830),
    .X(net224));
 sky130_fd_sc_hd__and2_2 c25 (.A(net943),
    .B(net941),
    .X(net0));
 sky130_fd_sc_hd__mux4_2 c250 (.A0(net997),
    .A1(net1046),
    .A2(net77),
    .A3(net1180),
    .S0(net187),
    .S1(net112),
    .X(net225));
 sky130_fd_sc_hd__mux4_2 c251 (.A0(net10),
    .A1(net1061),
    .A2(net85),
    .A3(net208),
    .S0(net983),
    .S1(net853),
    .X(net226));
 sky130_fd_sc_hd__mux4_1 c252 (.A0(net92),
    .A1(net105),
    .A2(net23),
    .A3(net1057),
    .S0(net847),
    .S1(clknet_1_0__leaf_net854),
    .X(net227));
 sky130_fd_sc_hd__mux4_1 c253 (.A0(net171),
    .A1(net92),
    .A2(net204),
    .A3(net209),
    .S0(clknet_1_0__leaf_net227),
    .S1(net1010),
    .X(net228));
 sky130_fd_sc_hd__mux4_1 c254 (.A0(net135),
    .A1(clknet_1_0__leaf_net227),
    .A2(net152),
    .A3(net776),
    .S0(net849),
    .S1(net853),
    .X(net229));
 sky130_fd_sc_hd__mux4_1 c255 (.A0(net1090),
    .A1(net992),
    .A2(clknet_1_0__leaf_net229),
    .A3(net75),
    .S0(net853),
    .S1(net857),
    .X(net230));
 sky130_fd_sc_hd__mux4_1 c256 (.A0(net209),
    .A1(clknet_1_0__leaf_net96),
    .A2(net135),
    .A3(net92),
    .S0(clknet_1_0__leaf_net227),
    .S1(net1037),
    .X(net958));
 sky130_fd_sc_hd__mux4_1 c257 (.A0(net1181),
    .A1(clknet_1_0__leaf_net96),
    .A2(net77),
    .A3(net983),
    .S0(clknet_1_0__leaf_net228),
    .S1(net1002),
    .X(net231));
 sky130_fd_sc_hd__mux4_1 c258 (.A0(net204),
    .A1(net152),
    .A2(clknet_1_1__leaf_net96),
    .A3(net162),
    .S0(net1182),
    .S1(net830),
    .X(net232));
 sky130_fd_sc_hd__mux4_1 c259 (.A0(net89),
    .A1(net85),
    .A2(net113),
    .A3(clknet_1_0__leaf_net227),
    .S0(clknet_1_0__leaf_net232),
    .S1(clknet_1_0__leaf_net855),
    .X(net233));
 sky130_fd_sc_hd__and2_2 c26 (.A(net1062),
    .B(net8),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c260 (.A0(net85),
    .A1(net209),
    .A2(clknet_1_1__leaf_net215),
    .A3(net104),
    .S0(clknet_1_0__leaf_net232),
    .S1(net861),
    .X(net234));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(net176),
    .A1(clknet_1_1__leaf_net215),
    .A2(net85),
    .A3(clknet_1_0__leaf_net232),
    .S1(net859),
    .X(net235));
 sky130_fd_sc_hd__mux4_1 c262 (.A0(clknet_1_1__leaf_net229),
    .A1(clknet_1_0__leaf_net958),
    .A2(net164),
    .A3(net85),
    .S0(net777),
    .S1(net864),
    .X(net236));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net983),
    .A1(net1092),
    .A2(clknet_1_1__leaf_net232),
    .A3(net1053),
    .S0(net864),
    .S1(net865),
    .X(net237));
 sky130_fd_sc_hd__and2_1 c264 (.A(net1057),
    .B(net122),
    .X(net238));
 sky130_fd_sc_hd__and2_2 c265 (.A(net1061),
    .B(net238),
    .X(net239));
 sky130_fd_sc_hd__and2_4 c266 (.A(net123),
    .B(net1044),
    .X(net240));
 sky130_fd_sc_hd__and2_2 c267 (.A(net1060),
    .B(net124),
    .X(net241));
 sky130_fd_sc_hd__and2_2 c268 (.A(net241),
    .B(net1026),
    .X(net242));
 sky130_fd_sc_hd__and2_1 c269 (.A(net951),
    .B(net114),
    .X(net243));
 sky130_fd_sc_hd__and2_2 c27 (.A(net945),
    .B(net1),
    .X(net2));
 sky130_fd_sc_hd__and2_1 c270 (.A(net930),
    .B(net114),
    .X(net244));
 sky130_fd_sc_hd__or4bb_4 c271 (.A(net949),
    .B(net243),
    .C_N(net1055),
    .D_N(net1020),
    .X(net245));
 sky130_fd_sc_hd__and2_2 c272 (.A(net243),
    .B(net113),
    .X(net246));
 sky130_fd_sc_hd__and2_2 c273 (.A(net238),
    .B(net244),
    .X(net247));
 sky130_fd_sc_hd__and2_4 c274 (.A(net1020),
    .B(net1044),
    .X(net248));
 sky130_fd_sc_hd__and2_4 c275 (.A(net244),
    .B(net1065),
    .X(net249));
 sky130_fd_sc_hd__and2_4 c276 (.A(net248),
    .B(net239),
    .X(net250));
 sky130_fd_sc_hd__a2111o_4 c277 (.A1(net113),
    .A2(net245),
    .B1(net249),
    .C1(net1013),
    .D1(net1126),
    .X(net251));
 sky130_fd_sc_hd__and2_1 c278 (.A(net107),
    .B(net1020),
    .X(net252));
 sky130_fd_sc_hd__or4bb_4 c279 (.A(net116),
    .B(net247),
    .C_N(net249),
    .D_N(net1020),
    .X(net962));
 sky130_fd_sc_hd__and2_4 c28 (.A(net1059),
    .B(net1),
    .X(net3));
 sky130_fd_sc_hd__a2111o_1 c280 (.A1(net249),
    .A2(net238),
    .B1(net933),
    .C1(net1024),
    .D1(net124),
    .X(net253));
 sky130_fd_sc_hd__or4bb_4 c281 (.A(net1021),
    .B(net252),
    .C_N(net962),
    .D_N(net1013),
    .X(net254));
 sky130_fd_sc_hd__mux4_2 c282 (.A0(net251),
    .A1(net254),
    .A2(net1013),
    .A3(net1126),
    .S0(net1020),
    .S1(net1047),
    .X(net255));
 sky130_fd_sc_hd__a2111o_1 c283 (.A1(net253),
    .A2(net123),
    .B1(net251),
    .C1(net1013),
    .D1(net255),
    .X(net256));
 sky130_fd_sc_hd__and2_2 c284 (.A(net252),
    .B(net253),
    .X(net257));
 sky130_fd_sc_hd__or4bb_4 c285 (.A(net256),
    .B(net1104),
    .C_N(net242),
    .D_N(net951),
    .X(net258));
 sky130_fd_sc_hd__and2_1 c286 (.A(net951),
    .B(net11),
    .X(net259));
 sky130_fd_sc_hd__and2_4 c287 (.A(net9),
    .B(net121),
    .X(net260));
 sky130_fd_sc_hd__or4bb_4 c288 (.A(net933),
    .B(net121),
    .C_N(net122),
    .D_N(net1025),
    .X(net261));
 sky130_fd_sc_hd__a2111o_4 c289 (.A1(net253),
    .A2(net146),
    .B1(net11),
    .C1(net943),
    .D1(net122),
    .X(net963));
 sky130_fd_sc_hd__and2_4 c29 (.A(net943),
    .B(net944),
    .X(net4));
 sky130_fd_sc_hd__and3_4 c290 (.A(net1062),
    .B(net261),
    .C(net1009),
    .X(net262));
 sky130_fd_sc_hd__and3_1 c291 (.A(net145),
    .B(net9),
    .C(net1022),
    .X(net263));
 sky130_fd_sc_hd__and3_2 c292 (.A(net8),
    .B(net125),
    .C(net1009),
    .X(net264));
 sky130_fd_sc_hd__a2111o_1 c293 (.A1(net11),
    .A2(net0),
    .B1(net264),
    .C1(net1016),
    .D1(net1013),
    .X(net265));
 sky130_fd_sc_hd__and3_1 c294 (.A(net1016),
    .B(net131),
    .C(net1100),
    .X(net266));
 sky130_fd_sc_hd__and3_2 c295 (.A(net265),
    .B(net261),
    .C(net260),
    .X(net267));
 sky130_fd_sc_hd__and3_2 c296 (.A(net129),
    .B(net146),
    .C(net261),
    .X(net268));
 sky130_fd_sc_hd__a2111o_1 c297 (.A1(net1064),
    .A2(net1040),
    .B1(net265),
    .C1(net128),
    .D1(net264),
    .X(net269));
 sky130_fd_sc_hd__a2111o_2 c298 (.A1(net264),
    .A2(net11),
    .B1(net269),
    .C1(net267),
    .D1(net1016),
    .X(net270));
 sky130_fd_sc_hd__and3_1 c299 (.A(net267),
    .B(net933),
    .C(net264),
    .X(net973));
 sky130_fd_sc_hd__and2_4 c30 (.A(net0),
    .B(net3),
    .X(net5));
 sky130_fd_sc_hd__or4bb_2 c300 (.A(net939),
    .B(net1104),
    .C_N(net267),
    .D_N(net998),
    .X(net271));
 sky130_fd_sc_hd__a2111o_4 c301 (.A1(net248),
    .A2(net962),
    .B1(net270),
    .C1(net998),
    .D1(net142),
    .X(net272));
 sky130_fd_sc_hd__mux4_2 c302 (.A0(net1100),
    .A1(net242),
    .A2(net268),
    .A3(net267),
    .S0(net1052),
    .S1(net939),
    .X(net273));
 sky130_fd_sc_hd__a2111o_1 c303 (.A1(net1038),
    .A2(net265),
    .B1(net270),
    .C1(net273),
    .D1(net998),
    .X(net274));
 sky130_fd_sc_hd__mux4_2 c304 (.A0(net274),
    .A1(net273),
    .A2(net963),
    .A3(net253),
    .S0(net242),
    .S1(net1025),
    .X(net275));
 sky130_fd_sc_hd__a2111o_2 c305 (.A1(net272),
    .A2(net274),
    .B1(net275),
    .C1(net273),
    .D1(net998),
    .X(net276));
 sky130_fd_sc_hd__a2111o_2 c306 (.A1(net146),
    .A2(net272),
    .B1(net276),
    .C1(net275),
    .D1(net1026),
    .X(net277));
 sky130_fd_sc_hd__mux4_2 c307 (.A0(net269),
    .A1(net272),
    .A2(net274),
    .A3(net271),
    .S0(net277),
    .S1(net275),
    .X(net278));
 sky130_fd_sc_hd__and3_1 c308 (.A(net154),
    .B(net163),
    .C(net1025),
    .X(net279));
 sky130_fd_sc_hd__a2111o_1 c309 (.A1(net267),
    .A2(net990),
    .B1(net1091),
    .C1(net278),
    .D1(net169),
    .X(net280));
 sky130_fd_sc_hd__and2_4 c31 (.A(net5),
    .B(net1022),
    .X(net6));
 sky130_fd_sc_hd__a2111o_2 c310 (.A1(net127),
    .A2(net985),
    .B1(net1016),
    .C1(net1127),
    .D1(net791),
    .X(net281));
 sky130_fd_sc_hd__and3_2 c311 (.A(net131),
    .B(net1022),
    .C(net990),
    .X(net282));
 sky130_fd_sc_hd__mux4_2 c312 (.A0(net1018),
    .A1(net1155),
    .A2(net1022),
    .A3(net990),
    .S0(net257),
    .S1(net1127),
    .X(net283));
 sky130_fd_sc_hd__and3_1 c313 (.A(net243),
    .B(net118),
    .C(net264),
    .X(net284));
 sky130_fd_sc_hd__and3_1 c314 (.A(net141),
    .B(net113),
    .C(net282),
    .X(net285));
 sky130_fd_sc_hd__and3_2 c315 (.A(net168),
    .B(net281),
    .C(net1060),
    .X(net286));
 sky130_fd_sc_hd__and3_1 c316 (.A(net137),
    .B(net277),
    .C(net1127),
    .X(net287));
 sky130_fd_sc_hd__and3_2 c317 (.A(net34),
    .B(net281),
    .C(net136),
    .X(net288));
 sky130_fd_sc_hd__and2_2 c318 (.A(net117),
    .B(net285),
    .X(net289));
 sky130_fd_sc_hd__and3_2 c319 (.A(net930),
    .B(net287),
    .C(net36),
    .X(net290));
 sky130_fd_sc_hd__and2_4 c32 (.A(net1022),
    .B(net8),
    .X(net7));
 sky130_fd_sc_hd__buf_1 c320 (.A(net791),
    .X(net291));
 sky130_fd_sc_hd__and3_1 c321 (.A(net284),
    .B(net267),
    .C(net285),
    .X(net292));
 sky130_fd_sc_hd__and3_2 c322 (.A(net19),
    .B(net998),
    .C(net159),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_1 c323 (.A(net791),
    .X(net294));
 sky130_fd_sc_hd__mux4_2 c324 (.A0(net292),
    .A1(net266),
    .A2(net288),
    .A3(net21),
    .S0(net951),
    .S1(net260),
    .X(net295));
 sky130_fd_sc_hd__and3_1 c325 (.A(net150),
    .B(net262),
    .C(net288),
    .X(net296));
 sky130_fd_sc_hd__mux4_2 c326 (.A0(net294),
    .A1(net293),
    .A2(net1007),
    .A3(net106),
    .S0(net284),
    .S1(net168),
    .X(net297));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(net282),
    .A1(net293),
    .A2(net19),
    .A3(net286),
    .S0(net290),
    .S1(net1104),
    .X(net298));
 sky130_fd_sc_hd__buf_1 c328 (.A(clknet_1_0__leaf_net798),
    .X(net299));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net299),
    .A1(net267),
    .A2(net294),
    .A3(net243),
    .S0(net290),
    .S1(net242),
    .X(net300));
 sky130_fd_sc_hd__and2_2 c33 (.A(net1055),
    .B(net1038),
    .X(net8));
 sky130_fd_sc_hd__or4bb_1 c330 (.A(net282),
    .B(net291),
    .C_N(net32),
    .D_N(net1030),
    .X(net301));
 sky130_fd_sc_hd__or4bb_1 c331 (.A(net278),
    .B(net1195),
    .C_N(net1155),
    .D_N(net1036),
    .X(net302));
 sky130_fd_sc_hd__a2111o_2 c332 (.A1(net1194),
    .A2(net156),
    .B1(net990),
    .C1(net939),
    .D1(net106),
    .X(net953));
 sky130_fd_sc_hd__a2111o_1 c333 (.A1(net138),
    .A2(net282),
    .B1(net273),
    .C1(net246),
    .D1(net982),
    .X(net303));
 sky130_fd_sc_hd__mux4_2 c334 (.A0(net21),
    .A1(net134),
    .A2(net155),
    .A3(net990),
    .S0(net1038),
    .S1(net997),
    .X(net304));
 sky130_fd_sc_hd__or4bb_2 c335 (.A(net301),
    .B(net178),
    .C_N(net989),
    .D_N(net145),
    .X(net305));
 sky130_fd_sc_hd__mux4_1 c336 (.A0(net254),
    .A1(net145),
    .A2(net987),
    .A3(net157),
    .S0(net296),
    .S1(net1036),
    .X(net306));
 sky130_fd_sc_hd__a2111o_1 c337 (.A1(net1051),
    .A2(net48),
    .B1(net990),
    .C1(net271),
    .D1(net1041),
    .X(net307));
 sky130_fd_sc_hd__a2111o_1 c338 (.A1(net271),
    .A2(net989),
    .B1(net939),
    .C1(net34),
    .D1(net1038),
    .X(net308));
 sky130_fd_sc_hd__a2111o_1 c339 (.A1(net302),
    .A2(net183),
    .B1(net141),
    .C1(net1096),
    .D1(clknet_1_0__leaf_net797),
    .X(net309));
 sky130_fd_sc_hd__and3_2 c34 (.A(net3),
    .B(net5),
    .C(net1062),
    .X(net9));
 sky130_fd_sc_hd__a2111o_1 c340 (.A1(net291),
    .A2(net41),
    .B1(net282),
    .C1(net175),
    .D1(net1030),
    .X(net310));
 sky130_fd_sc_hd__a2111o_1 c341 (.A1(net303),
    .A2(net290),
    .B1(net930),
    .C1(net987),
    .D1(net1030),
    .X(net311));
 sky130_fd_sc_hd__mux4_1 c342 (.A0(net7),
    .A1(net969),
    .A2(net153),
    .A3(net308),
    .S0(net1064),
    .S1(net310),
    .X(net312));
 sky130_fd_sc_hd__mux4_1 c343 (.A0(net32),
    .A1(net292),
    .A2(net28),
    .A3(net977),
    .S0(net308),
    .S1(net307),
    .X(net313));
 sky130_fd_sc_hd__mux4_1 c344 (.A0(net302),
    .A1(net257),
    .A2(net977),
    .A3(net1030),
    .S0(net1143),
    .S1(net1029),
    .X(net314));
 sky130_fd_sc_hd__mux4_1 c345 (.A0(net290),
    .A1(net939),
    .A2(net990),
    .A3(net1017),
    .S0(net842),
    .S1(net1029),
    .X(net315));
 sky130_fd_sc_hd__mux4_1 c346 (.A0(net191),
    .A1(net159),
    .A2(net977),
    .A3(net254),
    .S0(net1011),
    .S1(net1029),
    .X(net316));
 sky130_fd_sc_hd__mux4_1 c347 (.A0(net310),
    .A1(net56),
    .A2(net977),
    .A3(net1010),
    .S0(net138),
    .S1(net1029),
    .X(net317));
 sky130_fd_sc_hd__a2111o_1 c348 (.A1(net273),
    .A2(net1009),
    .B1(net977),
    .C1(net824),
    .D1(net1029),
    .X(net318));
 sky130_fd_sc_hd__mux4_1 c349 (.A0(net977),
    .A1(net6),
    .A2(net1082),
    .A3(net1198),
    .S0(net832),
    .S1(net1029),
    .X(net319));
 sky130_fd_sc_hd__or4bb_4 c35 (.A(net5),
    .B(net7),
    .C_N(net1047),
    .D_N(net6),
    .X(net10));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(net141),
    .A1(net291),
    .A2(net302),
    .A3(net977),
    .S0(net964),
    .S1(net832),
    .X(net320));
 sky130_fd_sc_hd__a2111o_1 c351 (.A1(net254),
    .A2(net803),
    .B1(net832),
    .C1(net842),
    .D1(net867),
    .X(net321));
 sky130_fd_sc_hd__a2111o_1 c352 (.A1(net70),
    .A2(net996),
    .B1(net207),
    .C1(net987),
    .D1(net1040),
    .X(net322));
 sky130_fd_sc_hd__a2111o_4 c353 (.A1(net261),
    .A2(net68),
    .B1(net207),
    .C1(net251),
    .D1(net851),
    .X(net323));
 sky130_fd_sc_hd__mux4_2 c354 (.A0(net257),
    .A1(net239),
    .A2(net6),
    .A3(net1059),
    .S0(net198),
    .S1(net1017),
    .X(net324));
 sky130_fd_sc_hd__mux4_2 c355 (.A0(net6),
    .A1(net930),
    .A2(net1042),
    .A3(net251),
    .S0(net1011),
    .S1(net842),
    .X(net325));
 sky130_fd_sc_hd__mux4_2 c356 (.A0(net134),
    .A1(net49),
    .A2(net282),
    .A3(net50),
    .S0(net1094),
    .S1(net1003),
    .X(net326));
 sky130_fd_sc_hd__mux4_2 c357 (.A0(net207),
    .A1(net67),
    .A2(net1085),
    .A3(net324),
    .S0(net930),
    .S1(net852),
    .X(net327));
 sky130_fd_sc_hd__a2111o_1 c358 (.A1(net325),
    .A2(net988),
    .B1(net207),
    .C1(net112),
    .D1(clknet_1_1__leaf_net797),
    .X(net328));
 sky130_fd_sc_hd__a2111o_1 c359 (.A1(net67),
    .A2(net996),
    .B1(net325),
    .C1(net1011),
    .D1(net73),
    .X(net329));
 sky130_fd_sc_hd__mux4_2 c36 (.A0(net1041),
    .A1(net10),
    .A2(net1038),
    .A3(net3),
    .S0(net943),
    .S1(net8),
    .X(net11));
 sky130_fd_sc_hd__mux4_1 c360 (.A0(net174),
    .A1(net945),
    .A2(net32),
    .A3(net1059),
    .S0(net1010),
    .S1(net65),
    .X(net330));
 sky130_fd_sc_hd__a2111o_1 c361 (.A1(net330),
    .A2(net239),
    .B1(net174),
    .C1(net1096),
    .D1(net322),
    .X(net331));
 sky130_fd_sc_hd__a2111o_1 c362 (.A1(net308),
    .A2(net32),
    .B1(net312),
    .C1(net41),
    .D1(net1036),
    .X(net332));
 sky130_fd_sc_hd__mux4_2 c363 (.A0(net331),
    .A1(net1159),
    .A2(net323),
    .A3(net1041),
    .S0(net1096),
    .S1(net1024),
    .X(net333));
 sky130_fd_sc_hd__mux4_1 c364 (.A0(net328),
    .A1(net1041),
    .A2(net977),
    .A3(net1036),
    .S0(net1054),
    .S1(net331),
    .X(net334));
 sky130_fd_sc_hd__a2111o_1 c365 (.A1(net329),
    .A2(net174),
    .B1(net1003),
    .C1(net51),
    .D1(net851),
    .X(net335));
 sky130_fd_sc_hd__mux4_1 c366 (.A0(net325),
    .A1(net144),
    .A2(net1004),
    .A3(net1018),
    .S0(net1061),
    .S1(net852),
    .X(net336));
 sky130_fd_sc_hd__a2111o_1 c367 (.A1(net336),
    .A2(net977),
    .B1(net1024),
    .C1(net1004),
    .D1(net200),
    .X(net337));
 sky130_fd_sc_hd__mux4_1 c368 (.A0(net277),
    .A1(net336),
    .A2(net987),
    .A3(net2),
    .S0(net70),
    .S1(clknet_1_1__leaf_net797),
    .X(net338));
 sky130_fd_sc_hd__a2111o_1 c369 (.A1(net335),
    .A2(net78),
    .B1(net325),
    .C1(net1011),
    .D1(net336),
    .X(net339));
 sky130_fd_sc_hd__and2_2 c37 (.A(net10),
    .B(net0),
    .X(net12));
 sky130_fd_sc_hd__a2111o_1 c370 (.A1(net112),
    .A2(net192),
    .B1(net1049),
    .C1(net838),
    .D1(net842),
    .X(net340));
 sky130_fd_sc_hd__a2111o_1 c371 (.A1(net340),
    .A2(net1049),
    .B1(net324),
    .C1(net115),
    .D1(net1031),
    .X(net341));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net1072),
    .A1(net340),
    .A2(net989),
    .A3(net32),
    .S0(net333),
    .S1(net838),
    .X(net342));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net340),
    .A1(net56),
    .A2(net1000),
    .A3(net325),
    .S0(net1007),
    .S1(net841),
    .X(net343));
 sky130_fd_sc_hd__mux4_1 c374 (.A0(clknet_1_1__leaf_net228),
    .A1(net1003),
    .A2(clknet_1_1__leaf_net96),
    .A3(net226),
    .S0(net1021),
    .S1(net1069),
    .X(net344));
 sky130_fd_sc_hd__mux4_1 c375 (.A0(net2),
    .A1(net1060),
    .A2(net323),
    .A3(clknet_1_1__leaf_net95),
    .S0(net982),
    .S1(net852),
    .X(net345));
 sky130_fd_sc_hd__mux4_1 c376 (.A0(clknet_1_1__leaf_net96),
    .A1(net326),
    .A2(net945),
    .A3(net162),
    .S0(clknet_1_0__leaf_net856),
    .S1(net860),
    .X(net346));
 sky130_fd_sc_hd__a2111o_1 c377 (.A1(net105),
    .A2(clknet_1_1__leaf_net346),
    .B1(net135),
    .C1(net970),
    .D1(net785),
    .X(net347));
 sky130_fd_sc_hd__mux4_1 c378 (.A0(net275),
    .A1(net105),
    .A2(net997),
    .A3(net1061),
    .S0(net828),
    .S1(net868),
    .X(net348));
 sky130_fd_sc_hd__mux4_1 c379 (.A0(net296),
    .A1(clknet_1_0__leaf_net227),
    .A2(clknet_1_0__leaf_net228),
    .A3(clknet_1_0__leaf_net95),
    .S0(net54),
    .S1(net864),
    .X(net349));
 sky130_fd_sc_hd__and3_4 c38 (.A(net6),
    .B(net943),
    .C(net10),
    .X(net13));
 sky130_fd_sc_hd__mux4_1 c380 (.A0(net226),
    .A1(net970),
    .A2(clknet_1_0__leaf_net222),
    .A3(net1010),
    .S0(net86),
    .S1(clknet_1_0__leaf_net232),
    .X(net350));
 sky130_fd_sc_hd__mux4_1 c381 (.A0(net54),
    .A1(net23),
    .A2(clknet_1_1__leaf_net95),
    .A3(net118),
    .S0(net975),
    .S1(net863),
    .X(net351));
 sky130_fd_sc_hd__mux4_1 c382 (.A0(net197),
    .A1(net982),
    .A2(net84),
    .A3(net135),
    .S0(clknet_1_1__leaf_net856),
    .S1(net868),
    .X(net352));
 sky130_fd_sc_hd__mux4_1 c383 (.A0(net50),
    .A1(net124),
    .A2(net246),
    .A3(net785),
    .S0(net817),
    .S1(net828),
    .X(net353));
 sky130_fd_sc_hd__mux4_1 c384 (.A0(net152),
    .A1(net75),
    .A2(net1073),
    .A3(net50),
    .S0(clknet_1_0__leaf_net346),
    .S1(net1059),
    .X(net354));
 sky130_fd_sc_hd__mux4_1 c385 (.A0(net49),
    .A1(clknet_1_1__leaf_net227),
    .A2(net225),
    .A3(net1070),
    .S0(clknet_1_1__leaf_net96),
    .S1(net853),
    .X(net355));
 sky130_fd_sc_hd__mux4_1 c386 (.A0(net86),
    .A1(net355),
    .A2(net92),
    .A3(net104),
    .S0(net226),
    .S1(clknet_1_0__leaf_net856),
    .X(net356));
 sky130_fd_sc_hd__mux4_1 c387 (.A0(net158),
    .A1(net982),
    .A2(net853),
    .A3(clknet_1_0__leaf_net855),
    .S0(net858),
    .S1(net864),
    .X(net357));
 sky130_fd_sc_hd__mux4_1 c388 (.A0(net56),
    .A1(net51),
    .A2(net86),
    .A3(net1198),
    .S0(net816),
    .S1(net965),
    .X(net358));
 sky130_fd_sc_hd__mux4_1 c389 (.A0(net6),
    .A1(net162),
    .A2(clknet_1_0__leaf_net222),
    .A3(clknet_1_1__leaf_net96),
    .S0(net817),
    .S1(net965),
    .X(net359));
 sky130_fd_sc_hd__and2_2 c39 (.A(net13),
    .B(net9),
    .X(net14));
 sky130_fd_sc_hd__mux4_1 c390 (.A0(clknet_1_1__leaf_net222),
    .A1(net338),
    .A2(net288),
    .A3(net325),
    .S0(net850),
    .S1(net870),
    .X(net957));
 sky130_fd_sc_hd__mux4_1 c391 (.A0(clknet_1_1__leaf_net95),
    .A1(net162),
    .A2(net785),
    .A3(net852),
    .S0(net864),
    .S1(net870),
    .X(net360));
 sky130_fd_sc_hd__mux4_1 c392 (.A0(net92),
    .A1(net322),
    .A2(net982),
    .A3(net1046),
    .S0(net869),
    .S1(net871),
    .X(net361));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net361),
    .A1(net1092),
    .A2(net982),
    .A3(net929),
    .S0(net858),
    .S1(net965),
    .X(net362));
 sky130_fd_sc_hd__mux4_1 c394 (.A0(net982),
    .A1(net75),
    .A2(net152),
    .A3(net964),
    .S0(net871),
    .S1(net965),
    .X(net363));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net359),
    .A1(net977),
    .A2(net363),
    .A3(clknet_1_0__leaf_net346),
    .S0(net1010),
    .S1(net965),
    .X(net364));
 sky130_fd_sc_hd__and2_2 c396 (.A(net1065),
    .B(net247),
    .X(net365));
 sky130_fd_sc_hd__and2_0 c397 (.A(net122),
    .B(net933),
    .X(net366));
 sky130_fd_sc_hd__and2_2 c398 (.A(net1055),
    .B(net241),
    .X(net367));
 sky130_fd_sc_hd__and3_1 c399 (.A(net108),
    .B(net366),
    .C(net123),
    .X(net368));
 sky130_fd_sc_hd__or4bb_4 c40 (.A(net944),
    .B(net14),
    .C_N(net6),
    .D_N(net8),
    .X(net15));
 sky130_fd_sc_hd__and2_1 c400 (.A(net368),
    .B(net121),
    .X(net369));
 sky130_fd_sc_hd__and2_0 c401 (.A(net252),
    .B(net366),
    .X(net370));
 sky130_fd_sc_hd__and2_2 c402 (.A(net949),
    .B(net107),
    .X(net371));
 sky130_fd_sc_hd__and2_4 c403 (.A(net258),
    .B(net252),
    .X(net372));
 sky130_fd_sc_hd__or4bb_4 c404 (.A(net119),
    .B(net372),
    .C_N(net251),
    .D_N(net962),
    .X(net373));
 sky130_fd_sc_hd__and3_2 c405 (.A(net117),
    .B(net370),
    .C(net1026),
    .X(net374));
 sky130_fd_sc_hd__and2_1 c406 (.A(net256),
    .B(net365),
    .X(net375));
 sky130_fd_sc_hd__and2_1 c407 (.A(net369),
    .B(net373),
    .X(net376));
 sky130_fd_sc_hd__and2_2 c408 (.A(net365),
    .B(net123),
    .X(net377));
 sky130_fd_sc_hd__a2111o_1 c409 (.A1(net373),
    .A2(net256),
    .B1(net368),
    .C1(net108),
    .D1(net1015),
    .X(net378));
 sky130_fd_sc_hd__mux4_2 c41 (.A0(net14),
    .A1(net13),
    .A2(net15),
    .A3(net944),
    .S0(net1059),
    .S1(net0),
    .X(net16));
 sky130_fd_sc_hd__a2111o_1 c410 (.A1(net1015),
    .A2(net369),
    .B1(net994),
    .C1(net1052),
    .D1(net121),
    .X(net379));
 sky130_fd_sc_hd__or4bb_4 c411 (.A(net121),
    .B(net256),
    .C_N(net371),
    .D_N(net994),
    .X(net380));
 sky130_fd_sc_hd__mux4_2 c412 (.A0(net238),
    .A1(net1015),
    .A2(net365),
    .A3(net994),
    .S0(net1065),
    .S1(net1005),
    .X(net381));
 sky130_fd_sc_hd__mux4_2 c413 (.A0(net380),
    .A1(net381),
    .A2(net1015),
    .A3(net365),
    .S0(net1005),
    .S1(net994),
    .X(net382));
 sky130_fd_sc_hd__or4bb_4 c414 (.A(net379),
    .B(net381),
    .C_N(net1015),
    .D_N(net994),
    .X(net383));
 sky130_fd_sc_hd__mux4_2 c415 (.A0(net372),
    .A1(net244),
    .A2(net383),
    .A3(net380),
    .S0(net365),
    .S1(net367),
    .X(net384));
 sky130_fd_sc_hd__mux4_2 c416 (.A0(net383),
    .A1(net382),
    .A2(net1008),
    .A3(net949),
    .S0(net1015),
    .S1(net1049),
    .X(net385));
 sky130_fd_sc_hd__mux4_2 c417 (.A0(net376),
    .A1(net384),
    .A2(net379),
    .A3(net1005),
    .S0(net365),
    .S1(net383),
    .X(net386));
 sky130_fd_sc_hd__and2_2 c418 (.A(net1060),
    .B(net128),
    .X(net387));
 sky130_fd_sc_hd__and3_1 c419 (.A(net121),
    .B(net269),
    .C(net1011),
    .X(net388));
 sky130_fd_sc_hd__and3_2 c42 (.A(net1052),
    .B(net1127),
    .C(net1055),
    .X(net17));
 sky130_fd_sc_hd__and3_1 c420 (.A(net380),
    .B(net371),
    .C(net1064),
    .X(net389));
 sky130_fd_sc_hd__a2111o_2 c421 (.A1(net265),
    .A2(net264),
    .B1(net270),
    .C1(net963),
    .D1(net254),
    .X(net390));
 sky130_fd_sc_hd__and3_1 c422 (.A(net1058),
    .B(net1065),
    .C(net1011),
    .X(net391));
 sky130_fd_sc_hd__mux4_2 c423 (.A0(net366),
    .A1(net270),
    .A2(net1009),
    .A3(net993),
    .S0(net1040),
    .S1(net1100),
    .X(net392));
 sky130_fd_sc_hd__and3_2 c424 (.A(net370),
    .B(net4),
    .C(net1112),
    .X(net393));
 sky130_fd_sc_hd__and2_2 c425 (.A(net274),
    .B(net1058),
    .X(net394));
 sky130_fd_sc_hd__and3_2 c426 (.A(net255),
    .B(net7),
    .C(net1131),
    .X(net395));
 sky130_fd_sc_hd__and3_2 c427 (.A(net128),
    .B(net268),
    .C(net1062),
    .X(net396));
 sky130_fd_sc_hd__and3_1 c428 (.A(net269),
    .B(net1018),
    .C(net1005),
    .X(net397));
 sky130_fd_sc_hd__and3_1 c429 (.A(net245),
    .B(net257),
    .C(net274),
    .X(net398));
 sky130_fd_sc_hd__and2_4 c43 (.A(net1065),
    .B(net928),
    .X(net18));
 sky130_fd_sc_hd__a2111o_2 c430 (.A1(net123),
    .A2(net370),
    .B1(net993),
    .C1(net1040),
    .D1(net398),
    .X(net399));
 sky130_fd_sc_hd__a2111o_4 c431 (.A1(net122),
    .A2(net1023),
    .B1(net1112),
    .C1(net1049),
    .D1(net984),
    .X(net400));
 sky130_fd_sc_hd__and3_1 c432 (.A(net397),
    .B(net392),
    .C(net7),
    .X(net401));
 sky130_fd_sc_hd__a2111o_2 c433 (.A1(net273),
    .A2(net122),
    .B1(net401),
    .C1(net1000),
    .D1(net0),
    .X(net402));
 sky130_fd_sc_hd__and3_1 c434 (.A(net7),
    .B(net398),
    .C(net393),
    .X(net403));
 sky130_fd_sc_hd__mux4_2 c435 (.A0(net257),
    .A1(net998),
    .A2(net1023),
    .A3(net1065),
    .S0(net394),
    .S1(net395),
    .X(net404));
 sky130_fd_sc_hd__a2111o_1 c436 (.A1(net403),
    .A2(net391),
    .B1(net398),
    .C1(net392),
    .D1(net1023),
    .X(net405));
 sky130_fd_sc_hd__a2111o_1 c437 (.A1(net1053),
    .A2(net1023),
    .B1(net404),
    .C1(net405),
    .D1(net1048),
    .X(net406));
 sky130_fd_sc_hd__a2111o_2 c438 (.A1(net404),
    .A2(net241),
    .B1(net367),
    .C1(net1016),
    .D1(net403),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net393),
    .A1(net407),
    .A2(net400),
    .A3(net1023),
    .S0(net401),
    .S1(net1041),
    .X(net408));
 sky130_fd_sc_hd__and3_2 c44 (.A(net1007),
    .B(net31),
    .C(net37),
    .X(net19));
 sky130_fd_sc_hd__and3_1 c440 (.A(net401),
    .B(net266),
    .C(net239),
    .X(net409));
 sky130_fd_sc_hd__or4bb_1 c441 (.A(net16),
    .B(net1021),
    .C_N(net791),
    .D_N(net814),
    .X(net410));
 sky130_fd_sc_hd__and3_1 c442 (.A(net369),
    .B(net389),
    .C(net386),
    .X(net411));
 sky130_fd_sc_hd__mux4_2 c443 (.A0(net410),
    .A1(net29),
    .A2(net377),
    .A3(net112),
    .S0(net151),
    .S1(net380),
    .X(net412));
 sky130_fd_sc_hd__mux4_1 c444 (.A0(net405),
    .A1(net1000),
    .A2(net159),
    .A3(net1055),
    .S0(net295),
    .S1(net40),
    .X(net413));
 sky130_fd_sc_hd__mux4_1 c445 (.A0(net389),
    .A1(net409),
    .A2(net29),
    .A3(net367),
    .S0(net401),
    .S1(net136),
    .X(net414));
 sky130_fd_sc_hd__or4bb_2 c446 (.A(net414),
    .B(net264),
    .C_N(net1023),
    .D_N(net412),
    .X(net415));
 sky130_fd_sc_hd__or4bb_1 c447 (.A(net130),
    .B(net1046),
    .C_N(net287),
    .D_N(net410),
    .X(net416));
 sky130_fd_sc_hd__sdfrbp_2 c448 (.CLK(clknet_4_2_0_clk),
    .D(net416),
    .RESET_B(net29),
    .SCD(net118),
    .SCE(net997),
    .Q(net418),
    .Q_N(net417));
 sky130_fd_sc_hd__or4bb_2 c449 (.A(net130),
    .B(net287),
    .C_N(net415),
    .D_N(net787),
    .X(net419));
 sky130_fd_sc_hd__a2111o_2 c45 (.A1(net29),
    .A2(net28),
    .B1(net26),
    .C1(net928),
    .D1(net5),
    .X(net20));
 sky130_fd_sc_hd__a2111o_1 c450 (.A1(net266),
    .A2(net239),
    .B1(net415),
    .C1(net406),
    .D1(net416),
    .X(net420));
 sky130_fd_sc_hd__and3_2 c451 (.A(net40),
    .B(net266),
    .C(net1025),
    .X(net421));
 sky130_fd_sc_hd__mux4_2 c452 (.A0(net264),
    .A1(net242),
    .A2(net985),
    .A3(net1005),
    .S0(net272),
    .S1(net292),
    .X(net422));
 sky130_fd_sc_hd__or4bb_4 c453 (.A(net998),
    .B(net400),
    .C_N(net421),
    .D_N(net787),
    .X(net423));
 sky130_fd_sc_hd__mux4_1 c454 (.A0(net409),
    .A1(net1166),
    .A2(net159),
    .A3(net981),
    .S0(net257),
    .S1(net395),
    .X(net424));
 sky130_fd_sc_hd__sdfbbn_1 c455 (.CLK_N(clknet_4_9_0_clk),
    .D(net424),
    .RESET_B(net418),
    .SCD(net981),
    .SCE(net111),
    .SET_B(net787),
    .Q(net426),
    .Q_N(net425));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(net287),
    .A1(net418),
    .A2(net389),
    .A3(net286),
    .S0(net981),
    .S1(net814),
    .X(net427));
 sky130_fd_sc_hd__or4bb_4 c457 (.A(net981),
    .B(net268),
    .C_N(net425),
    .D_N(net791),
    .X(net428));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(net411),
    .A1(net367),
    .A2(net258),
    .A3(net428),
    .S0(net281),
    .S1(net981),
    .X(net429));
 sky130_fd_sc_hd__and3_1 c459 (.A(net401),
    .B(net421),
    .C(net814),
    .X(net430));
 sky130_fd_sc_hd__mux4_2 c46 (.A0(net1),
    .A1(net36),
    .A2(net939),
    .A3(net15),
    .S0(net31),
    .S1(net1047),
    .X(net21));
 sky130_fd_sc_hd__mux4_2 c460 (.A0(net430),
    .A1(net986),
    .A2(net981),
    .A3(net156),
    .S0(net1026),
    .S1(net814),
    .X(net431));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net414),
    .A1(net431),
    .A2(net157),
    .A3(net23),
    .S0(net787),
    .S1(net814),
    .X(net432));
 sky130_fd_sc_hd__a2111o_1 c462 (.A1(net285),
    .A2(net49),
    .B1(net943),
    .C1(net1025),
    .D1(net997),
    .X(net433));
 sky130_fd_sc_hd__or4bb_1 c463 (.A(net33),
    .B(net995),
    .C_N(net417),
    .D_N(net1030),
    .X(net434));
 sky130_fd_sc_hd__mux4_2 c464 (.A0(net394),
    .A1(net112),
    .A2(net987),
    .A3(net1008),
    .S0(net1029),
    .S1(net867),
    .X(net435));
 sky130_fd_sc_hd__a2111o_1 c465 (.A1(net191),
    .A2(net162),
    .B1(net434),
    .C1(net155),
    .D1(net824),
    .X(net436));
 sky130_fd_sc_hd__a2111o_2 c466 (.A1(net305),
    .A2(net127),
    .B1(net7),
    .C1(net1024),
    .D1(net394),
    .X(net437));
 sky130_fd_sc_hd__a2111o_1 c467 (.A1(net1000),
    .A2(net305),
    .B1(net191),
    .C1(net107),
    .D1(net814),
    .X(net438));
 sky130_fd_sc_hd__a2111o_1 c468 (.A1(net1041),
    .A2(net1198),
    .B1(net976),
    .C1(net438),
    .D1(clknet_1_0__leaf_net797),
    .X(net439));
 sky130_fd_sc_hd__mux4_2 c469 (.A0(net943),
    .A1(net434),
    .A2(net371),
    .A3(net990),
    .S0(net1188),
    .S1(net127),
    .X(net440));
 sky130_fd_sc_hd__a2111o_4 c47 (.A1(net31),
    .A2(net39),
    .B1(net38),
    .C1(net1041),
    .D1(net30),
    .X(net22));
 sky130_fd_sc_hd__mux4_1 c470 (.A0(net25),
    .A1(net48),
    .A2(net157),
    .A3(net1062),
    .S0(net1049),
    .S1(net1031),
    .X(net441));
 sky130_fd_sc_hd__a2111o_1 c471 (.A1(net178),
    .A2(net153),
    .B1(net1040),
    .C1(net976),
    .D1(net139),
    .X(net442));
 sky130_fd_sc_hd__mux4_2 c472 (.A0(net441),
    .A1(net157),
    .A2(net371),
    .A3(net48),
    .S0(net1049),
    .S1(net35),
    .X(net443));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(net242),
    .A1(net1005),
    .A2(net976),
    .A3(net279),
    .S0(net380),
    .S1(net824),
    .X(net444));
 sky130_fd_sc_hd__a2111o_1 c474 (.A1(net1098),
    .A2(net1000),
    .B1(net305),
    .C1(net976),
    .D1(net1036),
    .X(net445));
 sky130_fd_sc_hd__a2111o_1 c475 (.A1(net995),
    .A2(net433),
    .B1(net48),
    .C1(net1051),
    .D1(net976),
    .X(net446));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(net380),
    .A1(net415),
    .A2(net987),
    .A3(net976),
    .S0(net386),
    .S1(net822),
    .X(net447));
 sky130_fd_sc_hd__sdfbbp_1 c477 (.CLK(clknet_4_2_0_clk),
    .D(net406),
    .RESET_B(net262),
    .SCD(net273),
    .SCE(net1064),
    .SET_B(net976),
    .Q(net449),
    .Q_N(net448));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(net45),
    .A1(net1046),
    .A2(net448),
    .A3(net417),
    .S0(net1116),
    .S1(net767),
    .X(net450));
 sky130_fd_sc_hd__sdfbbn_2 c479 (.CLK_N(clknet_4_3_0_clk),
    .D(net436),
    .RESET_B(net39),
    .SCD(net449),
    .SCE(net415),
    .SET_B(net440),
    .Q(net955),
    .Q_N(net451));
 sky130_fd_sc_hd__or4bb_4 c48 (.A(net9),
    .B(net35),
    .C_N(net38),
    .D_N(net1127),
    .X(net23));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net433),
    .A1(net415),
    .A2(net285),
    .A3(net45),
    .S0(net451),
    .S1(net1008),
    .X(net452));
 sky130_fd_sc_hd__mux4_2 c481 (.A0(net151),
    .A1(net976),
    .A2(net441),
    .A3(net435),
    .S0(net987),
    .S1(net1029),
    .X(net453));
 sky130_fd_sc_hd__mux4_2 c482 (.A0(net428),
    .A1(net451),
    .A2(net1009),
    .A3(net976),
    .S0(net1036),
    .S1(net829),
    .X(net454));
 sky130_fd_sc_hd__a2111o_1 c483 (.A1(net321),
    .A2(net273),
    .B1(net448),
    .C1(net804),
    .D1(net832),
    .X(net455));
 sky130_fd_sc_hd__mux4_1 c484 (.A0(net415),
    .A1(net1067),
    .A2(net987),
    .A3(net989),
    .S0(net986),
    .S1(net1031),
    .X(net456));
 sky130_fd_sc_hd__mux4_2 c485 (.A0(net1167),
    .A1(net1040),
    .A2(net449),
    .A3(net1049),
    .S0(net1036),
    .S1(net993),
    .X(net457));
 sky130_fd_sc_hd__mux4_1 c486 (.A0(net292),
    .A1(net1000),
    .A2(net993),
    .A3(net1066),
    .S0(net16),
    .S1(net1061),
    .X(net458));
 sky130_fd_sc_hd__mux4_2 c487 (.A0(net68),
    .A1(net81),
    .A2(net440),
    .A3(net1057),
    .S0(net989),
    .S1(net873),
    .X(net459));
 sky130_fd_sc_hd__mux4_2 c488 (.A0(net990),
    .A1(net124),
    .A2(net1066),
    .A3(net1061),
    .S0(net1116),
    .S1(net851),
    .X(net460));
 sky130_fd_sc_hd__mux4_1 c489 (.A0(net73),
    .A1(net79),
    .A2(net997),
    .A3(net933),
    .S0(net829),
    .S1(net852),
    .X(net461));
 sky130_fd_sc_hd__a2111o_1 c49 (.A1(net1064),
    .A2(net10),
    .B1(net34),
    .C1(net11),
    .D1(net21),
    .X(net24));
 sky130_fd_sc_hd__mux4_1 c490 (.A0(net987),
    .A1(net257),
    .A2(net260),
    .A3(net407),
    .S0(net35),
    .S1(net995),
    .X(net462));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(net449),
    .A1(net333),
    .A2(net1095),
    .A3(net407),
    .S0(clknet_1_0__leaf_net966),
    .S1(net852),
    .X(net463));
 sky130_fd_sc_hd__mux4_1 c492 (.A0(net262),
    .A1(net1159),
    .A2(net139),
    .A3(net1188),
    .S0(net1007),
    .S1(net823),
    .X(net464));
 sky130_fd_sc_hd__mux4_2 c493 (.A0(net239),
    .A1(net458),
    .A2(net326),
    .A3(net156),
    .S0(net459),
    .S1(net1004),
    .X(net465));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(net437),
    .A1(net212),
    .A2(net993),
    .A3(net760),
    .S0(net822),
    .S1(clknet_1_0__leaf_net966),
    .X(net466));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(net371),
    .A1(net333),
    .A2(net49),
    .A3(net465),
    .S0(net457),
    .S1(net933),
    .X(net467));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(net367),
    .A1(net438),
    .A2(net16),
    .A3(net115),
    .S0(net1040),
    .S1(clknet_1_0__leaf_net875),
    .X(net468));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net41),
    .A1(net465),
    .A2(net990),
    .A3(net1189),
    .S0(net760),
    .S1(clknet_1_0__leaf_net875),
    .X(net469));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(net456),
    .A1(net955),
    .A2(net452),
    .A3(net993),
    .S0(net1031),
    .S1(net851),
    .X(net470));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(net173),
    .A1(net1053),
    .A2(net440),
    .A3(net1060),
    .S0(net1031),
    .S1(clknet_1_1__leaf_net876),
    .X(net471));
 sky130_fd_sc_hd__a2111o_1 c50 (.A1(net928),
    .A2(net1064),
    .B1(net38),
    .C1(net32),
    .D1(net1046),
    .X(net25));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(net1051),
    .A1(net144),
    .A2(net324),
    .A3(net1031),
    .S0(net835),
    .S1(clknet_1_0__leaf_net876),
    .X(net472));
 sky130_fd_sc_hd__mux4_2 c501 (.A0(net212),
    .A1(net450),
    .A2(net987),
    .A3(net1031),
    .S0(clknet_1_0__leaf_net833),
    .S1(clknet_1_1__leaf_net876),
    .X(net473));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(net461),
    .A1(net452),
    .A2(net73),
    .A3(net459),
    .S0(clknet_1_0__leaf_net875),
    .S1(clknet_1_0__leaf_net876),
    .X(net474));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(net464),
    .A1(net988),
    .A2(net460),
    .A3(net304),
    .S0(net986),
    .S1(net836),
    .X(net475));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net386),
    .A1(net1102),
    .A2(net464),
    .A3(net304),
    .S0(net846),
    .S1(clknet_1_0__leaf_net876),
    .X(net476));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(net955),
    .A1(net456),
    .A2(net768),
    .A3(net823),
    .S0(net846),
    .S1(clknet_1_0__leaf_net875),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c506 (.A0(net164),
    .A1(net982),
    .A2(net327),
    .A3(net460),
    .S0(net421),
    .S1(net816),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c507 (.A0(net81),
    .A1(net23),
    .A2(net1040),
    .A3(clknet_1_1__leaf_net232),
    .S0(net84),
    .S1(net465),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c508 (.A0(net1025),
    .A1(net1024),
    .A2(net1096),
    .A3(net295),
    .S0(net353),
    .S1(net417),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c509 (.A0(net1073),
    .A1(net988),
    .A2(clknet_1_0__leaf_net352),
    .A3(net189),
    .S0(net863),
    .S1(clknet_1_1__leaf_net876),
    .X(net481));
 sky130_fd_sc_hd__and2_1 c51 (.A(net1051),
    .B(net38),
    .X(net26));
 sky130_fd_sc_hd__mux4_1 c510 (.A0(clknet_1_1__leaf_net232),
    .A1(clknet_1_0__leaf_net473),
    .A2(net976),
    .A3(net124),
    .S0(net1036),
    .S1(net865),
    .X(net482));
 sky130_fd_sc_hd__mux4_1 c511 (.A0(net1071),
    .A1(net999),
    .A2(clknet_1_1__leaf_net232),
    .A3(net288),
    .S0(net327),
    .S1(net853),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c512 (.A0(net407),
    .A1(net353),
    .A2(net437),
    .A3(net963),
    .S0(net1037),
    .S1(net260),
    .X(net484));
 sky130_fd_sc_hd__mux4_1 c513 (.A0(net358),
    .A1(net1061),
    .A2(net295),
    .A3(net831),
    .S0(net852),
    .S1(clknet_1_1__leaf_net876),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c514 (.A0(net348),
    .A1(net1049),
    .A2(net84),
    .A3(net963),
    .S0(net323),
    .S1(net878),
    .X(net486));
 sky130_fd_sc_hd__mux4_1 c515 (.A0(net437),
    .A1(net421),
    .A2(net288),
    .A3(net863),
    .S0(net877),
    .S1(net879),
    .X(net487));
 sky130_fd_sc_hd__mux4_1 c516 (.A0(net326),
    .A1(net1053),
    .A2(net407),
    .A3(net1054),
    .S0(net865),
    .S1(net872),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c517 (.A0(net162),
    .A1(net1036),
    .A2(net225),
    .A3(net295),
    .S0(net1004),
    .S1(net872),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c518 (.A0(net465),
    .A1(net363),
    .A2(net437),
    .A3(net81),
    .S0(net852),
    .S1(net879),
    .X(net490));
 sky130_fd_sc_hd__mux4_1 c519 (.A0(net295),
    .A1(clknet_1_1__leaf_net352),
    .A2(net190),
    .A3(net421),
    .S0(net1040),
    .S1(net883),
    .X(net491));
 sky130_fd_sc_hd__a2111o_4 c52 (.A1(net33),
    .A2(net24),
    .B1(net23),
    .C1(net1007),
    .D1(net1062),
    .X(net27));
 sky130_fd_sc_hd__mux4_1 c520 (.A0(clknet_1_1__leaf_net346),
    .A1(net988),
    .A2(clknet_1_1__leaf_net855),
    .A3(clknet_1_1__leaf_net874),
    .S0(net880),
    .S1(net883),
    .X(net492));
 sky130_fd_sc_hd__mux4_1 c521 (.A0(net327),
    .A1(net1036),
    .A2(clknet_1_1__leaf_net958),
    .A3(net853),
    .S0(net965),
    .S1(net883),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c522 (.A0(net84),
    .A1(net135),
    .A2(net460),
    .A3(net829),
    .S0(net862),
    .S1(net872),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c523 (.A0(net339),
    .A1(net113),
    .A2(net295),
    .A3(net995),
    .S0(clknet_1_0__leaf_net833),
    .S1(net880),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c524 (.A0(net1073),
    .A1(net118),
    .A2(net813),
    .A3(net831),
    .S0(net845),
    .S1(net864),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c525 (.A0(net288),
    .A1(net496),
    .A2(net1069),
    .A3(net1063),
    .S0(net864),
    .S1(net880),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c526 (.A0(net418),
    .A1(net17),
    .A2(net189),
    .A3(net81),
    .S0(net841),
    .S1(net845),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c527 (.A0(net421),
    .A1(net494),
    .A2(net81),
    .A3(net295),
    .S0(net869),
    .S1(net883),
    .X(net499));
 sky130_fd_sc_hd__and2_1 c528 (.A(net373),
    .B(net108),
    .X(net500));
 sky130_fd_sc_hd__and2_1 c529 (.A(net372),
    .B(net108),
    .X(net501));
 sky130_fd_sc_hd__and2_4 c53 (.A(net26),
    .B(net3),
    .X(net28));
 sky130_fd_sc_hd__and2_2 c530 (.A(net933),
    .B(net383),
    .X(net502));
 sky130_fd_sc_hd__and3_1 c531 (.A(net245),
    .B(net1064),
    .C(net502),
    .X(net503));
 sky130_fd_sc_hd__and3_4 c532 (.A(net247),
    .B(net1168),
    .C(net1021),
    .X(net504));
 sky130_fd_sc_hd__and2_0 c533 (.A(net379),
    .B(net116),
    .X(net505));
 sky130_fd_sc_hd__and2_1 c534 (.A(net505),
    .B(net245),
    .X(net506));
 sky130_fd_sc_hd__and3_4 c535 (.A(net984),
    .B(net384),
    .C(net1046),
    .X(net507));
 sky130_fd_sc_hd__and3_1 c536 (.A(net365),
    .B(net949),
    .C(net502),
    .X(net508));
 sky130_fd_sc_hd__and2_2 c537 (.A(net242),
    .B(net502),
    .X(net509));
 sky130_fd_sc_hd__and3_1 c538 (.A(net505),
    .B(net933),
    .C(net509),
    .X(net510));
 sky130_fd_sc_hd__a2111o_2 c539 (.A1(net248),
    .A2(net502),
    .B1(net1043),
    .C1(net365),
    .D1(net1049),
    .X(net511));
 sky130_fd_sc_hd__and3_2 c54 (.A(net1064),
    .B(net1038),
    .C(net5),
    .X(net29));
 sky130_fd_sc_hd__and2_1 c540 (.A(net381),
    .B(net510),
    .X(net512));
 sky130_fd_sc_hd__and2_2 c541 (.A(net368),
    .B(net504),
    .X(net513));
 sky130_fd_sc_hd__and3_1 c542 (.A(net376),
    .B(net507),
    .C(net1026),
    .X(net514));
 sky130_fd_sc_hd__sdfbbn_2 c543 (.CLK_N(clknet_4_8_0_clk),
    .D(net512),
    .RESET_B(net506),
    .SCD(net514),
    .SCE(net513),
    .SET_B(net502),
    .Q(net516),
    .Q_N(net515));
 sky130_fd_sc_hd__mux4_2 c544 (.A0(net510),
    .A1(net514),
    .A2(net504),
    .A3(net254),
    .S0(net502),
    .S1(net515),
    .X(net517));
 sky130_fd_sc_hd__a2111o_4 c545 (.A1(net511),
    .A2(net503),
    .B1(net1120),
    .C1(net1045),
    .D1(net1043),
    .X(net518));
 sky130_fd_sc_hd__mux4_1 c546 (.A0(net517),
    .A1(net518),
    .A2(net512),
    .A3(net1008),
    .S0(net970),
    .S1(net1118),
    .X(net519));
 sky130_fd_sc_hd__clkbuf_1 c547 (.A(net750),
    .X(net520));
 sky130_fd_sc_hd__and3_1 c548 (.A(net502),
    .B(net509),
    .C(net1112),
    .X(net521));
 sky130_fd_sc_hd__sdfbbp_1 c549 (.CLK(clknet_4_8_0_clk),
    .D(net506),
    .RESET_B(net376),
    .SCD(net521),
    .SCE(net368),
    .SET_B(net512),
    .Q(net523),
    .Q_N(net522));
 sky130_fd_sc_hd__and3_2 c55 (.A(net930),
    .B(net13),
    .C(net1047),
    .X(net30));
 sky130_fd_sc_hd__mux4_2 c550 (.A0(net388),
    .A1(net399),
    .A2(net276),
    .A3(net262),
    .S0(net1009),
    .S1(net500),
    .X(net524));
 sky130_fd_sc_hd__mux4_2 c551 (.A0(net514),
    .A1(net393),
    .A2(net518),
    .A3(net258),
    .S0(net254),
    .S1(net241),
    .X(net525));
 sky130_fd_sc_hd__mux4_2 c552 (.A0(net393),
    .A1(net391),
    .A2(net993),
    .A3(net507),
    .S0(net1093),
    .S1(net511),
    .X(net972));
 sky130_fd_sc_hd__mux4_1 c553 (.A0(net513),
    .A1(net1015),
    .A2(net1023),
    .A3(net107),
    .S0(net1132),
    .S1(net517),
    .X(net526));
 sky130_fd_sc_hd__mux4_2 c554 (.A0(net276),
    .A1(net1023),
    .A2(net984),
    .A3(net270),
    .S0(net515),
    .S1(net1055),
    .X(net527));
 sky130_fd_sc_hd__mux4_1 c555 (.A0(net1009),
    .A1(net136),
    .A2(net1015),
    .A3(net509),
    .S0(net1119),
    .S1(net979),
    .X(net528));
 sky130_fd_sc_hd__mux4_2 c556 (.A0(net244),
    .A1(net140),
    .A2(net979),
    .A3(net984),
    .S0(net522),
    .S1(net885),
    .X(net529));
 sky130_fd_sc_hd__mux4_1 c557 (.A0(net528),
    .A1(net147),
    .A2(net241),
    .A3(net1112),
    .S0(net1009),
    .S1(net527),
    .X(net530));
 sky130_fd_sc_hd__a2111o_1 c558 (.A1(net527),
    .A2(net393),
    .B1(net500),
    .C1(net529),
    .X(net531));
 sky130_fd_sc_hd__mux4_1 c559 (.A0(net398),
    .A1(net529),
    .A2(net525),
    .A3(net1098),
    .S0(net1016),
    .S1(net998),
    .X(net532));
 sky130_fd_sc_hd__and2_2 c56 (.A(net1061),
    .B(net29),
    .X(net31));
 sky130_fd_sc_hd__mux4_1 c560 (.A0(net528),
    .A1(net112),
    .A2(net518),
    .A3(net979),
    .S0(net754),
    .S1(net793),
    .X(net533));
 sky130_fd_sc_hd__mux4_2 c561 (.A0(net529),
    .A1(net527),
    .A2(net979),
    .A3(net1015),
    .S0(net754),
    .S1(net1028),
    .X(net534));
 sky130_fd_sc_hd__mux4_1 c562 (.A0(net500),
    .A1(net147),
    .A2(net516),
    .A3(net142),
    .S0(net793),
    .S1(net885),
    .X(net535));
 sky130_fd_sc_hd__mux4_2 c563 (.A0(net0),
    .A1(net1054),
    .A2(net1104),
    .A3(net793),
    .S0(net1028),
    .S1(net887),
    .X(net536));
 sky130_fd_sc_hd__mux4_1 c564 (.A0(net536),
    .A1(net503),
    .A2(net527),
    .A3(net1132),
    .S0(net276),
    .S1(net887),
    .X(net537));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net535),
    .A1(net527),
    .A2(net537),
    .A3(net518),
    .S0(net1028),
    .S1(net887),
    .X(net538));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(net108),
    .A1(net118),
    .A2(net536),
    .A3(net507),
    .S0(net1015),
    .S1(net1028),
    .X(net539));
 sky130_fd_sc_hd__mux4_1 c567 (.A0(net270),
    .A1(net524),
    .A2(net528),
    .A3(net393),
    .S0(net1132),
    .S1(net887),
    .X(net540));
 sky130_fd_sc_hd__mux4_2 c568 (.A0(net140),
    .A1(net1038),
    .A2(net262),
    .A3(net147),
    .S0(net1028),
    .S1(net889),
    .X(net541));
 sky130_fd_sc_hd__mux4_2 c569 (.A0(net539),
    .A1(net535),
    .A2(net536),
    .A3(net1098),
    .S0(net541),
    .S1(net754),
    .X(net542));
 sky130_fd_sc_hd__and2_2 c57 (.A(net7),
    .B(net951),
    .X(net32));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net536),
    .A1(net539),
    .A2(net248),
    .A3(net542),
    .S0(net754),
    .S1(net891),
    .X(net543));
 sky130_fd_sc_hd__mux4_1 c571 (.A0(net537),
    .A1(net539),
    .A2(net535),
    .A3(net517),
    .S0(net754),
    .S1(net892),
    .X(net544));
 sky130_fd_sc_hd__mux4_1 c572 (.A0(net412),
    .A1(net112),
    .A2(net1088),
    .A3(net513),
    .S0(net156),
    .S1(net890),
    .X(net545));
 sky130_fd_sc_hd__mux4_1 c573 (.A0(net29),
    .A1(net1183),
    .A2(net1064),
    .A3(net1046),
    .S0(net425),
    .S1(net1028),
    .X(net546));
 sky130_fd_sc_hd__mux4_1 c574 (.A0(net281),
    .A1(net541),
    .A2(net431),
    .A3(net515),
    .S0(net986),
    .S1(net887),
    .X(net547));
 sky130_fd_sc_hd__mux4_2 c575 (.A0(net399),
    .A1(net1060),
    .A2(net258),
    .A3(net240),
    .S0(net773),
    .S1(net885),
    .X(net548));
 sky130_fd_sc_hd__mux4_2 c576 (.A0(net39),
    .A1(net518),
    .A2(net377),
    .A3(net981),
    .S0(net515),
    .S1(net892),
    .X(net549));
 sky130_fd_sc_hd__mux4_1 c577 (.A0(net518),
    .A1(net545),
    .A2(net549),
    .A3(net431),
    .S0(net1063),
    .S1(net1028),
    .X(net550));
 sky130_fd_sc_hd__mux4_1 c578 (.A0(net136),
    .A1(net509),
    .A2(net281),
    .A3(net286),
    .S0(net283),
    .S1(net892),
    .X(net551));
 sky130_fd_sc_hd__mux4_1 c579 (.A0(net419),
    .A1(net422),
    .A2(net546),
    .A3(net4),
    .S0(net541),
    .S1(net143),
    .X(net552));
 sky130_fd_sc_hd__and2_4 c58 (.A(net30),
    .B(net941),
    .X(net33));
 sky130_fd_sc_hd__mux4_2 c580 (.A0(net162),
    .A1(net511),
    .A2(net39),
    .A3(net1018),
    .S0(net783),
    .S1(net1027),
    .X(net553));
 sky130_fd_sc_hd__mux4_2 c581 (.A0(net1052),
    .A1(net1008),
    .A2(net553),
    .A3(net993),
    .S0(net885),
    .S1(net1028),
    .X(net554));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(net399),
    .A1(net518),
    .A2(net515),
    .A3(net783),
    .S0(net888),
    .S1(net893),
    .X(net555));
 sky130_fd_sc_hd__mux4_1 c583 (.A0(net240),
    .A1(net553),
    .A2(net283),
    .A3(net981),
    .S0(net412),
    .S1(net825),
    .X(net556));
 sky130_fd_sc_hd__mux4_1 c584 (.A0(net286),
    .A1(net399),
    .A2(net1098),
    .A3(net981),
    .S0(net791),
    .S1(net893),
    .X(net557));
 sky130_fd_sc_hd__mux4_1 c585 (.A0(net120),
    .A1(net125),
    .A2(net419),
    .A3(net553),
    .S0(net554),
    .S1(net515),
    .X(net558));
 sky130_fd_sc_hd__mux4_1 c586 (.A0(net36),
    .A1(net549),
    .A2(net293),
    .A3(net1055),
    .S0(net1150),
    .S1(net1141),
    .X(net559));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(net556),
    .A1(net549),
    .A2(net541),
    .A3(net1016),
    .S0(net946),
    .S1(net773),
    .X(net560));
 sky130_fd_sc_hd__mux4_1 c588 (.A0(net503),
    .A1(net556),
    .A2(net258),
    .A3(net419),
    .S0(net518),
    .S1(net1046),
    .X(net561));
 sky130_fd_sc_hd__mux4_1 c589 (.A0(net147),
    .A1(net511),
    .A2(net159),
    .A3(net395),
    .S0(net894),
    .S1(clknet_1_0__leaf_net895),
    .X(net562));
 sky130_fd_sc_hd__and2_2 c59 (.A(net5),
    .B(net939),
    .X(net34));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(net1074),
    .A1(net1109),
    .A2(net136),
    .A3(net986),
    .S0(net773),
    .S1(clknet_1_0__leaf_net895),
    .X(net563));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(net545),
    .A1(net293),
    .A2(net39),
    .A3(net1051),
    .S0(net979),
    .S1(net773),
    .X(net564));
 sky130_fd_sc_hd__mux4_1 c592 (.A0(net555),
    .A1(net503),
    .A2(clknet_1_0__leaf_net563),
    .A3(net515),
    .S0(net839),
    .S1(clknet_1_0__leaf_net895),
    .X(net565));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(net150),
    .A1(net1023),
    .A2(net811),
    .A3(net825),
    .S0(net839),
    .S1(net893),
    .X(net566));
 sky130_fd_sc_hd__mux4_2 c594 (.A0(net142),
    .A1(net435),
    .A2(net1124),
    .A3(net867),
    .S0(net1027),
    .S1(net894),
    .X(net567));
 sky130_fd_sc_hd__mux4_2 c595 (.A0(net144),
    .A1(net399),
    .A2(net804),
    .A3(net824),
    .S0(net873),
    .S1(net889),
    .X(net568));
 sky130_fd_sc_hd__mux4_2 c596 (.A0(net307),
    .A1(net567),
    .A2(net1009),
    .A3(net1194),
    .S0(net811),
    .S1(net893),
    .X(net569));
 sky130_fd_sc_hd__mux4_1 c597 (.A0(net392),
    .A1(net938),
    .A2(net283),
    .A3(net513),
    .S0(net1011),
    .S1(net1130),
    .X(net570));
 sky130_fd_sc_hd__mux4_1 c598 (.A0(net377),
    .A1(net1163),
    .A2(net1130),
    .A3(net1087),
    .S0(net175),
    .S1(net839),
    .X(net571));
 sky130_fd_sc_hd__mux4_1 c599 (.A0(net509),
    .A1(net254),
    .A2(net549),
    .A3(net568),
    .S0(net832),
    .S1(net891),
    .X(net572));
 sky130_fd_sc_hd__and2_4 c60 (.A(net34),
    .B(net30),
    .X(net35));
 sky130_fd_sc_hd__mux4_2 c600 (.A0(net157),
    .A1(net1101),
    .A2(net567),
    .A3(net1098),
    .S0(net509),
    .S1(net892),
    .X(net573));
 sky130_fd_sc_hd__mux4_1 c601 (.A0(net549),
    .A1(net1008),
    .A2(net573),
    .A3(net307),
    .S0(net144),
    .S1(net893),
    .X(net574));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(net431),
    .A1(net1024),
    .A2(net569),
    .A3(net455),
    .S0(net814),
    .S1(clknet_1_0__leaf_net897),
    .X(net575));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(net183),
    .A1(net48),
    .A2(net259),
    .A3(net554),
    .S0(net513),
    .S1(net1027),
    .X(net576));
 sky130_fd_sc_hd__mux4_2 c604 (.A0(net48),
    .A1(net504),
    .A2(net455),
    .A3(net33),
    .S0(net47),
    .S1(net867),
    .X(net577));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net175),
    .A1(net27),
    .A2(net431),
    .A3(net1039),
    .S0(net885),
    .S1(clknet_1_0__leaf_net897),
    .X(net578));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net1184),
    .A1(net1017),
    .A2(net573),
    .A3(net435),
    .S0(net241),
    .S1(net803),
    .X(net579));
 sky130_fd_sc_hd__mux4_2 c607 (.A0(net567),
    .A1(net175),
    .A2(net451),
    .A3(net39),
    .S0(net806),
    .S1(net1029),
    .X(net580));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net509),
    .A1(net1039),
    .A2(net803),
    .A3(net824),
    .S0(net1027),
    .S1(net900),
    .X(net581));
 sky130_fd_sc_hd__mux4_1 c609 (.A0(net155),
    .A1(net159),
    .A2(net48),
    .A3(net1005),
    .S0(net573),
    .S1(net899),
    .X(net582));
 sky130_fd_sc_hd__and3_4 c61 (.A(net939),
    .B(net31),
    .C(net1022),
    .X(net36));
 sky130_fd_sc_hd__mux4_1 c610 (.A0(net241),
    .A1(net513),
    .A2(net142),
    .A3(net581),
    .S0(net567),
    .S1(net898),
    .X(net583));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net112),
    .A1(net573),
    .A2(net1124),
    .A3(net509),
    .S0(net577),
    .S1(clknet_1_0__leaf_net874),
    .X(net584));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(net283),
    .A1(net262),
    .A2(net1009),
    .A3(net567),
    .S0(net890),
    .S1(net904),
    .X(net585));
 sky130_fd_sc_hd__mux4_2 c613 (.A0(net455),
    .A1(net35),
    .A2(net392),
    .A3(net581),
    .S0(net175),
    .S1(net806),
    .X(net586));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(net581),
    .A1(net577),
    .A2(net549),
    .A3(net395),
    .S0(net1163),
    .S1(net443),
    .X(net587));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net583),
    .A1(net577),
    .A2(net1097),
    .A3(net803),
    .S0(net1141),
    .S1(clknet_1_0__leaf_net896),
    .X(net588));
 sky130_fd_sc_hd__mux4_1 c616 (.A0(net585),
    .A1(net111),
    .A2(net1129),
    .A3(net1051),
    .S0(net200),
    .S1(net988),
    .X(net589));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(net1014),
    .A1(net1106),
    .A2(net200),
    .A3(net324),
    .S0(net806),
    .S1(net893),
    .X(net590));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(net1056),
    .A1(net28),
    .A2(net585),
    .A3(net1061),
    .S0(net1053),
    .S1(net1136),
    .X(net591));
 sky130_fd_sc_hd__mux4_2 c619 (.A0(net79),
    .A1(net107),
    .A2(net1053),
    .A3(net323),
    .S0(net851),
    .S1(net888),
    .X(net592));
 sky130_fd_sc_hd__and2_2 c62 (.A(net9),
    .B(net30),
    .X(net37));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net592),
    .A1(net144),
    .A2(clknet_1_0__leaf_net471),
    .A3(net1063),
    .S0(net541),
    .S1(net443),
    .X(net593));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(net156),
    .A1(net1026),
    .A2(net374),
    .A3(net1007),
    .S0(net592),
    .S1(net516),
    .X(net594));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(net1086),
    .A1(net590),
    .A2(net190),
    .A3(net142),
    .S0(net982),
    .S1(net885),
    .X(net595));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(net993),
    .A1(net142),
    .A2(net1190),
    .A3(net65),
    .S0(net1129),
    .S1(net894),
    .X(net596));
 sky130_fd_sc_hd__mux4_1 c624 (.A0(net472),
    .A1(net1195),
    .A2(net190),
    .A3(net993),
    .S0(net132),
    .S1(net988),
    .X(net597));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net27),
    .A1(clknet_1_1__leaf_net597),
    .A2(net323),
    .A3(net1018),
    .S0(net1056),
    .S1(net1136),
    .X(net598));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net198),
    .A1(net541),
    .A2(net592),
    .A3(net262),
    .S0(net459),
    .S1(clknet_1_1__leaf_net897),
    .X(net967));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(net1049),
    .A1(net61),
    .A2(net569),
    .A3(net995),
    .S0(net836),
    .S1(net893),
    .X(net599));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(clknet_1_0__leaf_net597),
    .A1(net161),
    .A2(net190),
    .A3(net1103),
    .S0(net516),
    .S1(net804),
    .X(net600));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(net933),
    .A1(net116),
    .A2(net988),
    .A3(net460),
    .S0(net968),
    .S1(net905),
    .X(net601));
 sky130_fd_sc_hd__and2_2 c63 (.A(net943),
    .B(net30),
    .X(net38));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net1058),
    .A1(net66),
    .A2(net592),
    .A3(net988),
    .S0(net1086),
    .S1(clknet_1_0__leaf_net874),
    .X(net602));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net601),
    .A1(net1007),
    .A2(net516),
    .A3(net189),
    .S0(net788),
    .S1(net906),
    .X(net603));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net78),
    .A1(net986),
    .A2(net1129),
    .A3(net603),
    .S0(net440),
    .S1(net806),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(net603),
    .A1(net35),
    .A2(clknet_1_0__leaf_net593),
    .A3(net1107),
    .S0(net390),
    .S1(net844),
    .X(net605));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net260),
    .A1(net516),
    .A2(net16),
    .A3(net116),
    .S0(net786),
    .S1(net906),
    .X(net606));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net569),
    .A1(net28),
    .A2(net260),
    .A3(clknet_1_0__leaf_net967),
    .S0(clknet_1_1__leaf_net874),
    .S1(net902),
    .X(net607));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net65),
    .A1(net606),
    .A2(net200),
    .A3(net779),
    .S0(net905),
    .S1(net907),
    .X(net961));
 sky130_fd_sc_hd__mux4_2 c637 (.A0(net440),
    .A1(net65),
    .A2(net144),
    .A3(net841),
    .S0(net885),
    .S1(net907),
    .X(net608));
 sky130_fd_sc_hd__and2_4 c64 (.A(net1046),
    .B(net34),
    .X(net39));
 sky130_fd_sc_hd__mux4_1 c643 (.A0(net457),
    .A1(net1054),
    .A2(net947),
    .A3(net246),
    .S0(clknet_1_1__leaf_net833),
    .S1(net873),
    .X(net609));
 sky130_fd_sc_hd__mux4_1 c644 (.A0(net459),
    .A1(net478),
    .A2(net516),
    .A3(net850),
    .S0(net889),
    .S1(net907),
    .X(net610));
 sky130_fd_sc_hd__mux4_1 c645 (.A0(net1053),
    .A1(net486),
    .A2(net821),
    .A3(net835),
    .S0(net873),
    .S1(clknet_1_0__leaf_net896),
    .X(net611));
 sky130_fd_sc_hd__mux4_1 c646 (.A0(net1050),
    .A1(net1089),
    .A2(net988),
    .A3(net160),
    .S0(net841),
    .S1(net844),
    .X(net612));
 sky130_fd_sc_hd__mux4_1 c647 (.A0(net357),
    .A1(net1061),
    .A2(net611),
    .A3(net1097),
    .S0(net516),
    .S1(net839),
    .X(net613));
 sky130_fd_sc_hd__mux4_1 c648 (.A0(net260),
    .A1(net1004),
    .A2(net820),
    .A3(net850),
    .S0(net884),
    .S1(clknet_1_1__leaf_net896),
    .X(net614));
 sky130_fd_sc_hd__mux4_1 c649 (.A0(net142),
    .A1(net594),
    .A2(clknet_1_1__leaf_net227),
    .A3(net995),
    .S0(net881),
    .S1(net884),
    .X(net615));
 sky130_fd_sc_hd__and3_2 c65 (.A(net20),
    .B(net26),
    .C(net19),
    .X(net40));
 sky130_fd_sc_hd__mux4_1 c650 (.A0(net460),
    .A1(net541),
    .A2(net498),
    .A3(net1004),
    .S0(net828),
    .S1(net965),
    .X(net974));
 sky130_fd_sc_hd__mux4_1 c651 (.A0(net192),
    .A1(net516),
    .A2(net974),
    .A3(net1151),
    .S0(net873),
    .S1(net1142),
    .X(net616));
 sky130_fd_sc_hd__mux4_1 c652 (.A0(clknet_1_1__leaf_net471),
    .A1(net190),
    .A2(clknet_1_1__leaf_net563),
    .A3(net956),
    .S0(net1190),
    .S1(net882),
    .X(net617));
 sky130_fd_sc_hd__mux4_1 c653 (.A0(net931),
    .A1(net609),
    .A2(net982),
    .A3(net260),
    .S0(net807),
    .S1(net860),
    .X(net618));
 sky130_fd_sc_hd__mux4_1 c654 (.A0(net617),
    .A1(net486),
    .A2(net618),
    .A3(net132),
    .S0(net862),
    .S1(net891),
    .X(net619));
 sky130_fd_sc_hd__mux4_2 c655 (.A0(clknet_1_1__leaf_net473),
    .A1(net942),
    .A2(net1189),
    .A3(net995),
    .S0(net997),
    .S1(net849),
    .X(net620));
 sky130_fd_sc_hd__mux4_1 c656 (.A0(net497),
    .A1(net118),
    .A2(net323),
    .A3(net612),
    .S0(net827),
    .S1(net965),
    .X(net621));
 sky130_fd_sc_hd__mux4_1 c657 (.A0(net225),
    .A1(net1050),
    .A2(net821),
    .A3(net827),
    .S0(clknet_1_1__leaf_net874),
    .S1(net907),
    .X(net622));
 sky130_fd_sc_hd__mux4_1 c658 (.A0(net160),
    .A1(net614),
    .A2(net1014),
    .A3(clknet_1_0__leaf_net622),
    .S0(net190),
    .S1(net903),
    .X(net623));
 sky130_fd_sc_hd__mux4_1 c659 (.A0(net566),
    .A1(net112),
    .A2(clknet_1_1__leaf_net622),
    .A3(net778),
    .S0(clknet_1_0__leaf_net795),
    .S1(net837),
    .X(net624));
 sky130_fd_sc_hd__mux4_2 c66 (.A0(net59),
    .A1(net60),
    .A2(net55),
    .A3(net996),
    .S0(net46),
    .S1(net1034),
    .X(net969));
 sky130_fd_sc_hd__buf_1 c660 (.A(net762),
    .X(net625));
 sky130_fd_sc_hd__and3_1 c661 (.A(net1046),
    .B(net523),
    .C(net625),
    .X(net626));
 sky130_fd_sc_hd__and2_1 c662 (.A(net1169),
    .B(net626),
    .X(net627));
 sky130_fd_sc_hd__and3_1 c663 (.A(net125),
    .B(net1075),
    .C(net627),
    .X(net628));
 sky130_fd_sc_hd__or4bb_1 c664 (.A(net1056),
    .B(net1168),
    .C_N(net970),
    .D_N(net1054),
    .X(net629));
 sky130_fd_sc_hd__or4bb_1 c665 (.A(net629),
    .B(net1100),
    .C_N(net240),
    .D_N(net1006),
    .X(net630));
 sky130_fd_sc_hd__or4bb_4 c666 (.A(net1076),
    .B(net1008),
    .C_N(net1005),
    .D_N(net628),
    .X(net960));
 sky130_fd_sc_hd__mux4_1 c667 (.A0(net970),
    .A1(net376),
    .A2(net960),
    .A3(net628),
    .S0(net629),
    .S1(net1005),
    .X(net631));
 sky130_fd_sc_hd__or4bb_1 c668 (.A(net949),
    .B(net521),
    .C_N(net1065),
    .D_N(net630),
    .X(net632));
 sky130_fd_sc_hd__and3_2 c669 (.A(net626),
    .B(net629),
    .C(net508),
    .X(net633));
 sky130_fd_sc_hd__and2_2 c67 (.A(net38),
    .B(net35),
    .X(net41));
 sky130_fd_sc_hd__and2_0 c670 (.A(net521),
    .B(net626),
    .X(net634));
 sky130_fd_sc_hd__clkbuf_1 c671 (.A(net762),
    .X(net635));
 sky130_fd_sc_hd__sdfbbn_1 c672 (.CLK_N(clknet_4_10_0_clk),
    .D(net1052),
    .RESET_B(net960),
    .SCD(net1170),
    .SCE(net634),
    .SET_B(net762),
    .Q(net637),
    .Q_N(net636));
 sky130_fd_sc_hd__and2_2 c673 (.A(net637),
    .B(net762),
    .X(net638));
 sky130_fd_sc_hd__clkbuf_4 c674 (.A(net750),
    .X(net954));
 sky130_fd_sc_hd__sdfbbn_2 c675 (.CLK_N(clknet_4_10_0_clk),
    .D(net520),
    .RESET_B(net1144),
    .SCD(net954),
    .SCE(net632),
    .SET_B(net1021),
    .Q(net640),
    .Q_N(net639));
 sky130_fd_sc_hd__and2_0 c676 (.A(net1051),
    .B(net954),
    .X(net641));
 sky130_fd_sc_hd__or4bb_1 c677 (.A(net635),
    .B(net640),
    .C_N(net630),
    .D_N(net636),
    .X(net642));
 sky130_fd_sc_hd__and2_2 c678 (.A(net641),
    .B(net949),
    .X(net643));
 sky130_fd_sc_hd__mux4_1 c679 (.A0(net634),
    .A1(net637),
    .A2(net949),
    .A3(net954),
    .S0(net633),
    .S1(net641),
    .X(net644));
 sky130_fd_sc_hd__and2_0 c68 (.A(net1064),
    .B(net941),
    .X(net42));
 sky130_fd_sc_hd__mux4_1 c680 (.A0(net642),
    .A1(net643),
    .A2(net639),
    .A3(net1021),
    .S0(net1122),
    .S1(net908),
    .X(net645));
 sky130_fd_sc_hd__mux4_2 c681 (.A0(net1065),
    .A1(net643),
    .A2(net640),
    .A3(net508),
    .S0(net970),
    .S1(net910),
    .X(net646));
 sky130_fd_sc_hd__mux4_1 c682 (.A0(net627),
    .A1(net517),
    .A2(net1121),
    .A3(net1019),
    .S0(net1012),
    .S1(net963),
    .X(net647));
 sky130_fd_sc_hd__mux4_1 c683 (.A0(net402),
    .A1(net1052),
    .A2(net524),
    .A3(net1065),
    .S0(net908),
    .S1(net1149),
    .X(net648));
 sky130_fd_sc_hd__mux4_2 c684 (.A0(net396),
    .A1(net523),
    .A2(net639),
    .A3(net1100),
    .S0(net942),
    .S1(net16),
    .X(net649));
 sky130_fd_sc_hd__mux4_2 c685 (.A0(net625),
    .A1(net638),
    .A2(net1006),
    .A3(net524),
    .S0(net1121),
    .S1(net1045),
    .X(net650));
 sky130_fd_sc_hd__mux4_1 c686 (.A0(net501),
    .A1(net524),
    .A2(net1008),
    .A3(net649),
    .S0(net1123),
    .S1(net1065),
    .X(net651));
 sky130_fd_sc_hd__mux4_2 c687 (.A0(net523),
    .A1(net1006),
    .A2(net636),
    .A3(net648),
    .S0(net761),
    .S1(net792),
    .X(net652));
 sky130_fd_sc_hd__mux4_1 c688 (.A0(net648),
    .A1(net1023),
    .A2(net272),
    .A3(net542),
    .S0(net1039),
    .S1(net1138),
    .X(net653));
 sky130_fd_sc_hd__mux4_2 c689 (.A0(net1121),
    .A1(net643),
    .A2(net1021),
    .A3(net508),
    .S0(net751),
    .S1(net792),
    .X(net654));
 sky130_fd_sc_hd__and3_1 c69 (.A(net1059),
    .B(net945),
    .C(net1032),
    .X(net43));
 sky130_fd_sc_hd__mux4_2 c690 (.A0(net16),
    .A1(net963),
    .A2(net627),
    .A3(net639),
    .S0(net522),
    .S1(net396),
    .X(net655));
 sky130_fd_sc_hd__mux4_1 c691 (.A0(net542),
    .A1(net4),
    .A2(net1006),
    .A3(net978),
    .S0(net522),
    .S1(net761),
    .X(net656));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(net508),
    .A1(net937),
    .A2(net978),
    .A3(net633),
    .S0(net1008),
    .S1(net1153),
    .X(net657));
 sky130_fd_sc_hd__mux4_1 c693 (.A0(net525),
    .A1(net387),
    .A2(net1053),
    .A3(net1016),
    .S0(net761),
    .S1(net912),
    .X(net658));
 sky130_fd_sc_hd__mux4_2 c694 (.A0(net391),
    .A1(net1052),
    .A2(net627),
    .A3(net978),
    .S0(net396),
    .S1(net1097),
    .X(net659));
 sky130_fd_sc_hd__mux4_1 c695 (.A0(net524),
    .A1(net978),
    .A2(net504),
    .A3(net625),
    .S0(net792),
    .S1(net909),
    .X(net660));
 sky130_fd_sc_hd__mux4_1 c696 (.A0(net628),
    .A1(net640),
    .A2(net657),
    .A3(net954),
    .S0(net1006),
    .S1(net978),
    .X(net661));
 sky130_fd_sc_hd__mux4_1 c697 (.A0(net937),
    .A1(net132),
    .A2(net1132),
    .A3(net638),
    .S0(net649),
    .S1(net911),
    .X(net662));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(net525),
    .A1(net662),
    .A2(net636),
    .A3(net978),
    .S0(net751),
    .S1(net826),
    .X(net663));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(net657),
    .A1(net978),
    .A2(net1132),
    .A3(net1137),
    .S0(net1152),
    .S1(net1148),
    .X(net664));
 sky130_fd_sc_hd__and3_4 c70 (.A(net1022),
    .B(net20),
    .C(net1032),
    .X(net956));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net652),
    .A1(net523),
    .A2(net627),
    .A3(net1052),
    .S0(net636),
    .S1(net912),
    .X(net665));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(net662),
    .A1(net501),
    .A2(net249),
    .A3(net1012),
    .S0(net781),
    .S1(net912),
    .X(net666));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net660),
    .A1(net659),
    .A2(net1012),
    .A3(net1056),
    .S0(net978),
    .S1(net826),
    .X(net667));
 sky130_fd_sc_hd__mux4_2 c703 (.A0(net998),
    .A1(net508),
    .A2(net794),
    .A3(net826),
    .S0(net886),
    .S1(net913),
    .X(net668));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net387),
    .A1(net978),
    .A2(net289),
    .A3(net161),
    .S0(net143),
    .S1(net963),
    .X(net669));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(net23),
    .A1(net646),
    .A2(net1016),
    .A3(net668),
    .S0(net649),
    .S1(net801),
    .X(net670));
 sky130_fd_sc_hd__mux4_1 c706 (.A0(net426),
    .A1(net1043),
    .A2(net143),
    .A3(net639),
    .S0(net1014),
    .S1(net293),
    .X(net671));
 sky130_fd_sc_hd__mux4_1 c707 (.A0(net143),
    .A1(net954),
    .A2(net387),
    .A3(net761),
    .S0(net839),
    .S1(net1138),
    .X(net672));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(net40),
    .A1(net1056),
    .A2(net638),
    .A3(net107),
    .S0(net794),
    .S1(net913),
    .X(net673));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(net402),
    .A1(net659),
    .A2(net297),
    .A3(net998),
    .S0(net554),
    .S1(net801),
    .X(net674));
 sky130_fd_sc_hd__or4bb_4 c71 (.A(net15),
    .B(net43),
    .C_N(net33),
    .D_N(net1032),
    .X(net44));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net546),
    .A1(net1052),
    .A2(net542),
    .A3(net1135),
    .S0(net553),
    .S1(net825),
    .X(net675));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net143),
    .A1(net659),
    .A2(net548),
    .A3(net1134),
    .S0(net504),
    .S1(net1028),
    .X(net676));
 sky130_fd_sc_hd__mux4_2 c712 (.A0(net289),
    .A1(net1025),
    .A2(net1078),
    .A3(net638),
    .S0(net1133),
    .S1(net1054),
    .X(net677));
 sky130_fd_sc_hd__mux4_1 c713 (.A0(net637),
    .A1(net553),
    .A2(net649),
    .A3(net646),
    .S0(net668),
    .S1(net913),
    .X(net678));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(net40),
    .A1(net33),
    .A2(net504),
    .A3(net297),
    .S0(net1053),
    .S1(net801),
    .X(net679));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net646),
    .A1(net669),
    .A2(net637),
    .A3(net1006),
    .S0(net794),
    .S1(clknet_1_1__leaf_net895),
    .X(net680));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net638),
    .A1(net402),
    .A2(net297),
    .A3(net652),
    .S0(net932),
    .S1(net554),
    .X(net681));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net946),
    .A1(net16),
    .A2(net1081),
    .A3(net677),
    .S0(net794),
    .S1(clknet_1_1__leaf_net895),
    .X(net682));
 sky130_fd_sc_hd__mux4_2 c718 (.A0(net293),
    .A1(net671),
    .A2(net426),
    .A3(net1016),
    .S0(net1079),
    .S1(net892),
    .X(net683));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net677),
    .A1(net542),
    .A2(net1008),
    .A3(net825),
    .S0(net908),
    .S1(net915),
    .X(net684));
 sky130_fd_sc_hd__and2_2 c72 (.A(net1032),
    .B(net14),
    .X(net45));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net1080),
    .A1(net1063),
    .A2(net934),
    .A3(clknet_1_1__leaf_net895),
    .S0(net915),
    .S1(clknet_1_0__leaf_net916),
    .X(net685));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net422),
    .A1(net678),
    .A2(net677),
    .A3(net554),
    .S0(net978),
    .S1(net1028),
    .X(net686));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net1077),
    .A1(net650),
    .A2(net954),
    .A3(net794),
    .S0(net915),
    .S1(clknet_1_0__leaf_net917),
    .X(net687));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net297),
    .A1(net293),
    .A2(net651),
    .A3(net289),
    .S0(net40),
    .S1(net886),
    .X(net688));
 sky130_fd_sc_hd__mux4_2 c724 (.A0(net143),
    .A1(net981),
    .A2(net402),
    .A3(net1021),
    .S0(net908),
    .S1(net914),
    .X(net689));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net651),
    .A1(net643),
    .A2(net668),
    .A3(net554),
    .S0(net826),
    .S1(clknet_1_0__leaf_net917),
    .X(net690));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net633),
    .A1(net1039),
    .A2(net1054),
    .A3(net580),
    .S0(net668),
    .S1(net249),
    .X(net691));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net1125),
    .A1(net249),
    .A2(net633),
    .A3(net673),
    .S0(clknet_1_0__leaf_net562),
    .S1(net16),
    .X(net692));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net685),
    .A1(net955),
    .A2(net580),
    .A3(net633),
    .S0(net780),
    .S1(net1029),
    .X(net693));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(net395),
    .A1(net167),
    .A2(net568),
    .A3(net670),
    .S0(net655),
    .S1(net999),
    .X(net694));
 sky130_fd_sc_hd__a2111o_4 c73 (.A1(net45),
    .A2(net44),
    .B1(net996),
    .C1(net1032),
    .D1(net15),
    .X(net46));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net650),
    .A1(net542),
    .A2(net44),
    .A3(net249),
    .S0(net948),
    .S1(net826),
    .X(net695));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net553),
    .A1(clknet_1_1__leaf_net562),
    .A2(net1198),
    .A3(net272),
    .S0(net1012),
    .S1(net904),
    .X(net696));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(net687),
    .A1(net652),
    .A2(net36),
    .A3(net120),
    .S0(net677),
    .S1(clknet_1_1__leaf_net918),
    .X(net697));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net504),
    .A1(net47),
    .A2(net970),
    .A3(net247),
    .S0(net1101),
    .S1(net920),
    .X(net698));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(net698),
    .A1(net167),
    .A2(net247),
    .A3(net802),
    .S0(net904),
    .S1(clknet_1_0__leaf_net918),
    .X(net699));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net698),
    .A1(net999),
    .A2(net650),
    .A3(net839),
    .S0(net913),
    .S1(net914),
    .X(net700));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(net44),
    .A1(net677),
    .A2(net542),
    .A3(net1019),
    .S0(net784),
    .S1(net802),
    .X(net701));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net580),
    .A1(net1014),
    .A2(net33),
    .A3(net443),
    .S0(net901),
    .S1(net923),
    .X(net702));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net700),
    .A1(net249),
    .A2(net952),
    .A3(net954),
    .S0(net914),
    .S1(net925),
    .X(net703));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(net1005),
    .A1(net1021),
    .A2(net1039),
    .A3(net568),
    .S0(net810),
    .S1(net925),
    .X(net704));
 sky130_fd_sc_hd__and3_2 c74 (.A(net31),
    .B(net944),
    .C(net1032),
    .X(net47));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(net670),
    .A1(net633),
    .A2(net810),
    .A3(net1146),
    .S0(net899),
    .S1(clknet_1_0__leaf_net916),
    .X(net705));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(net672),
    .A1(net554),
    .A2(net960),
    .A3(net36),
    .S0(net919),
    .S1(net921),
    .X(net706));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(net659),
    .A1(net272),
    .A2(net132),
    .A3(clknet_1_0__leaf_net834),
    .S0(net901),
    .S1(net924),
    .X(net707));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(net683),
    .A1(net700),
    .A2(net1012),
    .A3(net794),
    .S0(net840),
    .S1(net892),
    .X(net708));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(net553),
    .A1(net956),
    .A2(net633),
    .A3(clknet_1_0__leaf_net834),
    .S0(net843),
    .S1(net925),
    .X(net709));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(net696),
    .A1(net41),
    .A2(net504),
    .A3(net120),
    .S0(net892),
    .S1(net913),
    .X(net710));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net153),
    .A1(net683),
    .A2(net827),
    .A3(clknet_1_1__leaf_net834),
    .S0(net840),
    .S1(net866),
    .X(net711));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(net33),
    .A1(net780),
    .A2(net827),
    .A3(net840),
    .S0(clknet_1_1__leaf_net916),
    .S1(net971),
    .X(net712));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net272),
    .A1(net41),
    .A2(net689),
    .A3(net435),
    .S0(net840),
    .S1(clknet_1_1__leaf_net875),
    .X(net713));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net643),
    .A1(net435),
    .A2(net586),
    .A3(clknet_1_0__leaf_net709),
    .S0(net788),
    .S1(net832),
    .X(net714));
 sky130_fd_sc_hd__and3_2 c75 (.A(net43),
    .B(net3),
    .C(net1032),
    .X(net48));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(net4),
    .A1(clknet_1_1__leaf_net593),
    .A2(net963),
    .A3(net1019),
    .S0(net23),
    .S1(net744),
    .X(net715));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net1040),
    .A1(net36),
    .A2(net443),
    .A3(net652),
    .S0(net1017),
    .S1(net374),
    .X(net716));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net161),
    .A1(net247),
    .A2(net699),
    .A3(net1063),
    .S0(net608),
    .S1(net61),
    .X(net717));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net548),
    .A1(net1056),
    .A2(net608),
    .A3(net586),
    .S0(clknet_1_1__leaf_net834),
    .S1(clknet_1_1__leaf_net875),
    .X(net718));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net324),
    .A1(net1108),
    .A2(net988),
    .A3(net1019),
    .S0(net920),
    .S1(net922),
    .X(net719));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(clknet_1_0__leaf_net712),
    .A1(net1043),
    .A2(net649),
    .A3(net954),
    .S0(net443),
    .S1(net1019),
    .X(net720));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net655),
    .A1(net28),
    .A2(net548),
    .A3(net784),
    .S0(clknet_1_1__leaf_net966),
    .S1(net924),
    .X(net721));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net374),
    .A1(net1017),
    .A2(net606),
    .A3(net161),
    .S0(net1056),
    .S1(net649),
    .X(net722));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net936),
    .A1(net1045),
    .A2(clknet_1_1__leaf_net720),
    .A3(net960),
    .S0(clknet_1_1__leaf_net795),
    .S1(net905),
    .X(net723));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net586),
    .A1(net655),
    .A2(clknet_1_0__leaf_net720),
    .A3(net805),
    .S0(net808),
    .S1(net926),
    .X(net724));
 sky130_fd_sc_hd__or4bb_4 c76 (.A(net1007),
    .B(net47),
    .C_N(net46),
    .D_N(net1033),
    .X(net49));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net1021),
    .A1(net689),
    .A2(net568),
    .A3(net324),
    .S0(net829),
    .S1(net1145),
    .X(net725));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net61),
    .A1(net704),
    .A2(net28),
    .A3(net1017),
    .S0(net837),
    .S1(net927),
    .X(net726));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net200),
    .A1(net692),
    .A2(net722),
    .A3(net1024),
    .S0(clknet_1_1__leaf_net712),
    .S1(net743),
    .X(net727));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(net1019),
    .A1(net946),
    .A2(net719),
    .A3(net586),
    .S0(net1115),
    .S1(net1140),
    .X(net728));
 sky130_fd_sc_hd__mux4_1 c764 (.A0(net673),
    .A1(net668),
    .A2(clknet_1_1__leaf_net709),
    .A3(net28),
    .S0(net324),
    .S1(net818),
    .X(net729));
 sky130_fd_sc_hd__mux4_1 c765 (.A0(clknet_1_1__leaf_net721),
    .A1(net1108),
    .A2(net786),
    .A3(clknet_1_1__leaf_net875),
    .S0(net905),
    .S1(clknet_1_1__leaf_net917),
    .X(net730));
 sky130_fd_sc_hd__mux4_1 c766 (.A0(net324),
    .A1(net819),
    .A2(net826),
    .A3(net843),
    .S0(clknet_1_1__leaf_net916),
    .S1(net971),
    .X(net731));
 sky130_fd_sc_hd__mux4_1 c767 (.A0(net652),
    .A1(net726),
    .A2(clknet_1_1__leaf_net731),
    .A3(net324),
    .S0(net813),
    .S1(clknet_1_1__leaf_net916),
    .X(net732));
 sky130_fd_sc_hd__mux4_1 c768 (.A0(net640),
    .A1(net568),
    .A2(net947),
    .A3(clknet_1_0__leaf_net731),
    .S0(net802),
    .S1(net805),
    .X(net733));
 sky130_fd_sc_hd__mux4_1 c769 (.A0(net41),
    .A1(net733),
    .A2(clknet_1_0__leaf_net721),
    .A3(net568),
    .S0(net804),
    .S1(clknet_1_1__leaf_net833),
    .X(net734));
 sky130_fd_sc_hd__and3_2 c77 (.A(net47),
    .B(net35),
    .C(net1032),
    .X(net50));
 sky130_fd_sc_hd__and3_2 c78 (.A(net39),
    .B(net43),
    .C(net1032),
    .X(net51));
 sky130_fd_sc_hd__a2111o_1 c79 (.A1(net26),
    .A2(net996),
    .B1(net31),
    .C1(net23),
    .D1(net1032),
    .X(net52));
 sky130_fd_sc_hd__or4bb_2 c80 (.A(net19),
    .B(net21),
    .C_N(net48),
    .D_N(net1033),
    .X(net53));
 sky130_fd_sc_hd__a2111o_2 c81 (.A1(net1010),
    .A2(net46),
    .B1(net52),
    .C1(net1034),
    .D1(net996),
    .X(net54));
 sky130_fd_sc_hd__and3_2 c82 (.A(net53),
    .B(net45),
    .C(net50),
    .X(net55));
 sky130_fd_sc_hd__or4bb_4 c83 (.A(net1058),
    .B(net55),
    .C_N(net44),
    .D_N(net1035),
    .X(net56));
 sky130_fd_sc_hd__mux4_2 c84 (.A0(net44),
    .A1(net1011),
    .A2(net53),
    .A3(net1060),
    .S0(net46),
    .S1(net55),
    .X(net57));
 sky130_fd_sc_hd__mux4_2 c85 (.A0(net57),
    .A1(net52),
    .A2(net45),
    .A3(net1034),
    .S0(net1010),
    .S1(net1055),
    .X(net58));
 sky130_fd_sc_hd__a2111o_2 c86 (.A1(net56),
    .A2(net58),
    .B1(net31),
    .C1(net1033),
    .D1(net1048),
    .X(net59));
 sky130_fd_sc_hd__mux4_2 c87 (.A0(net1010),
    .A1(net54),
    .A2(net52),
    .A3(net55),
    .S0(net59),
    .S1(net1034),
    .X(net60));
 sky130_fd_sc_hd__and2_2 c88 (.A(net16),
    .B(net46),
    .X(net61));
 sky130_fd_sc_hd__and2_0 c89 (.A(net1062),
    .B(net22),
    .X(net62));
 sky130_fd_sc_hd__and3_1 c90 (.A(net37),
    .B(net1033),
    .C(net996),
    .X(net63));
 sky130_fd_sc_hd__a2111o_1 c91 (.A1(net1011),
    .A2(net22),
    .B1(net991),
    .C1(net1034),
    .D1(net1001),
    .X(net64));
 sky130_fd_sc_hd__and2_2 c92 (.A(net1003),
    .B(net23),
    .X(net65));
 sky130_fd_sc_hd__and3_1 c93 (.A(net30),
    .B(net996),
    .C(net1001),
    .X(net66));
 sky130_fd_sc_hd__and2_1 c94 (.A(net1048),
    .B(net56),
    .X(net67));
 sky130_fd_sc_hd__and2_2 c95 (.A(net22),
    .B(net61),
    .X(net68));
 sky130_fd_sc_hd__and3_1 c96 (.A(net1110),
    .B(net68),
    .C(net1001),
    .X(net69));
 sky130_fd_sc_hd__and3_1 c97 (.A(net32),
    .B(net54),
    .C(net991),
    .X(net70));
 sky130_fd_sc_hd__and3_1 c98 (.A(net64),
    .B(net13),
    .C(net1001),
    .X(net71));
 sky130_fd_sc_hd__mux4_1 c99 (.A0(net1111),
    .A1(net6),
    .A2(net69),
    .A3(net991),
    .S0(net61),
    .S1(net1001),
    .X(net72));
 sky130_fd_sc_hd__a2111o_1 merge790 (.A1(net127),
    .A2(net8),
    .B1(net286),
    .C1(net289),
    .D1(net268),
    .X(net735));
 sky130_fd_sc_hd__a2111o_1 merge791 (.A1(net632),
    .A2(net625),
    .B1(net517),
    .C1(net520),
    .D1(net522),
    .X(net736));
 sky130_fd_sc_hd__mux4_1 merge792 (.A0(net515),
    .A1(net512),
    .A2(net365),
    .A3(net630),
    .S0(net632),
    .S1(net1139),
    .X(net737));
 sky130_fd_sc_hd__mux4_1 merge793 (.A0(net1180),
    .A1(net72),
    .A2(net89),
    .A3(net169),
    .S0(net278),
    .S1(net23),
    .X(net738));
 sky130_fd_sc_hd__and2_0 merge794 (.A(net695),
    .B(net703),
    .X(net739));
 sky130_fd_sc_hd__and2_0 merge795 (.A(net734),
    .B(net713),
    .X(net740));
 sky130_fd_sc_hd__and2_0 merge796 (.A(net332),
    .B(net334),
    .X(net741));
 sky130_fd_sc_hd__and2_0 merge797 (.A(net195),
    .B(net203),
    .X(net742));
 sky130_fd_sc_hd__dfrbp_1 merge798 (.CLK(clknet_4_12_0_clk),
    .D(net589),
    .RESET_B(net591),
    .Q(net744),
    .Q_N(net743));
 sky130_fd_sc_hd__and2_0 merge799 (.A(net574),
    .B(net575),
    .X(net745));
 sky130_fd_sc_hd__and2_0 merge800 (.A(net551),
    .B(net565),
    .X(net746));
 sky130_fd_sc_hd__and2_0 merge801 (.A(net610),
    .B(net613),
    .X(net747));
 sky130_fd_sc_hd__and2_0 merge802 (.A(net217),
    .B(net224),
    .X(net748));
 sky130_fd_sc_hd__and2_0 merge803 (.A(net309),
    .B(net315),
    .X(net749));
 sky130_fd_sc_hd__dfrbp_1 merge804 (.CLK(clknet_4_8_0_clk),
    .D(net519),
    .RESET_B(net737),
    .Q(net751),
    .Q_N(net750));
 sky130_fd_sc_hd__and2_0 merge805 (.A(net679),
    .B(net681),
    .X(net752));
 sky130_fd_sc_hd__and2_0 merge806 (.A(net439),
    .B(net442),
    .X(net753));
 sky130_fd_sc_hd__dfrtn_1 merge807 (.CLK_N(clknet_4_8_0_clk),
    .D(net530),
    .Q(net531));
 sky130_fd_sc_hd__and2_0 merge808 (.A(net345),
    .B(net350),
    .X(net755));
 sky130_fd_sc_hd__and2_0 merge809 (.A(net480),
    .B(net481),
    .X(net756));
 sky130_fd_sc_hd__and2_0 merge810 (.A(net186),
    .B(net185),
    .X(net757));
 sky130_fd_sc_hd__and2_0 merge811 (.A(net413),
    .B(net427),
    .X(net758));
 sky130_fd_sc_hd__and2_0 merge812 (.A(net280),
    .B(net735),
    .X(net759));
 sky130_fd_sc_hd__dfrtp_1 merge813 (.CLK(clknet_4_3_0_clk),
    .D(net462),
    .RESET_B(net463),
    .Q(net760));
 sky130_fd_sc_hd__dfrtp_2 merge814 (.CLK(clknet_4_10_0_clk),
    .D(net647),
    .RESET_B(net653),
    .Q(net761));
 sky130_fd_sc_hd__dfrtp_1 merge815 (.CLK(clknet_4_10_0_clk),
    .D(net736),
    .RESET_B(net631),
    .Q(net762));
 sky130_fd_sc_hd__dfsbp_1 merge816 (.CLK(clknet_4_4_0_clk),
    .D(net93),
    .Q(net101),
    .Q_N(net763));
 sky130_fd_sc_hd__and2_0 merge817 (.A(net454),
    .B(net447),
    .X(net765));
 sky130_fd_sc_hd__and2_0 merge818 (.A(net319),
    .B(net587),
    .X(net766));
 sky130_fd_sc_hd__dfsbp_1 merge819 (.CLK(clknet_4_3_0_clk),
    .D(net476),
    .SET_B(net445),
    .Q(net768),
    .Q_N(net767));
 sky130_fd_sc_hd__and2_0 merge820 (.A(net364),
    .B(net362),
    .X(net769));
 sky130_fd_sc_hd__and2_0 merge821 (.A(net690),
    .B(net682),
    .X(net770));
 sky130_fd_sc_hd__and2_0 merge822 (.A(net688),
    .B(net770),
    .X(net771));
 sky130_fd_sc_hd__and2_0 merge823 (.A(net337),
    .B(net605),
    .X(net772));
 sky130_fd_sc_hd__dfstp_1 merge824 (.CLK(clknet_4_9_0_clk),
    .D(net547),
    .SET_B(net559),
    .Q(net773));
 sky130_fd_sc_hd__and2_1 merge825 (.A(net343),
    .B(net499),
    .X(net774));
 sky130_fd_sc_hd__dfstp_1 merge826 (.CLK(clknet_4_13_0_clk),
    .D(net595),
    .SET_B(net624),
    .Q(net968));
 sky130_fd_sc_hd__dfstp_1 merge827 (.CLK(clknet_4_0_0_clk),
    .D(net188),
    .SET_B(net757),
    .Q(net775));
 sky130_fd_sc_hd__dlrbn_1 merge828 (.GATE_N(clknet_4_5_0_clk),
    .RESET_B(net748),
    .Q(net235),
    .Q_N(net776));
 sky130_fd_sc_hd__dlrbn_1 merge829 (.D(net604),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net623),
    .Q(net779),
    .Q_N(net778));
 sky130_fd_sc_hd__dlrbp_1 merge830 (.D(net661),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net752),
    .Q(net781),
    .Q_N(net780));
 sky130_fd_sc_hd__and2_0 merge831 (.A(net468),
    .B(net484),
    .X(net782));
 sky130_fd_sc_hd__dlrbp_1 merge832 (.D(net739),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net552),
    .Q(net784),
    .Q_N(net783));
 sky130_fd_sc_hd__dlrtn_1 merge833 (.D(net237),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net755),
    .Q(net785));
 sky130_fd_sc_hd__dlrtn_1 merge834 (.D(net729),
    .GATE_N(clknet_4_14_0_clk),
    .RESET_B(net598),
    .Q(net786));
 sky130_fd_sc_hd__dlrtn_2 merge835 (.D(net774),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net205),
    .Q(net975));
 sky130_fd_sc_hd__dlrtp_1 merge836 (.D(net420),
    .GATE(clknet_4_2_0_clk),
    .RESET_B(net758),
    .Q(net787));
 sky130_fd_sc_hd__dlrtp_1 merge837 (.D(net600),
    .GATE(clknet_4_14_0_clk),
    .RESET_B(net740),
    .Q(net788));
 sky130_fd_sc_hd__and2_0 merge838 (.A(net469),
    .B(net621),
    .X(net789));
 sky130_fd_sc_hd__and2_0 merge839 (.A(net474),
    .B(net477),
    .X(net790));
 sky130_fd_sc_hd__dlrtp_2 merge840 (.D(net759),
    .GATE(clknet_4_0_0_clk),
    .RESET_B(net298),
    .Q(net791));
 sky130_fd_sc_hd__edfxbp_1 merge841 (.CLK(clknet_4_8_0_clk),
    .D(net532),
    .DE(net544),
    .Q(net793),
    .Q_N(net792));
 sky130_fd_sc_hd__edfxtp_1 merge842 (.CLK(clknet_4_10_0_clk),
    .D(net667),
    .DE(net666),
    .Q(net794));
 sky130_fd_sc_hd__sdlclkp_1 merge843 (.CLK(clknet_4_15_0_clk),
    .GATE(net716),
    .SCE(net619),
    .GCLK(net795));
 sky130_fd_sc_hd__and2_0 merge844 (.A(net599),
    .B(net732),
    .X(net796));
 sky130_fd_sc_hd__sdlclkp_2 merge845 (.CLK(clknet_4_0_0_clk),
    .GATE(net306),
    .SCE(net311),
    .GCLK(net797));
 sky130_fd_sc_hd__sdlclkp_4 merge846 (.CLK(clknet_4_4_0_clk),
    .GATE(net214),
    .SCE(net738),
    .GCLK(net798));
 sky130_fd_sc_hd__dfrbp_1 merge847 (.CLK(clknet_4_1_0_clk),
    .D(net211),
    .RESET_B(net742),
    .Q(net800),
    .Q_N(net799));
 sky130_fd_sc_hd__dfrbp_2 merge848 (.CLK(clknet_4_10_0_clk),
    .D(net665),
    .RESET_B(net664),
    .Q(net802),
    .Q_N(net801));
 sky130_fd_sc_hd__dfrtn_1 merge849 (.CLK_N(clknet_4_12_0_clk),
    .D(net576),
    .RESET_B(net766),
    .Q(net803));
 sky130_fd_sc_hd__dfrtp_2 merge850 (.CLK(clknet_4_15_0_clk),
    .D(net796),
    .RESET_B(net453),
    .Q(net804));
 sky130_fd_sc_hd__dfrtp_1 merge851 (.CLK(clknet_4_15_0_clk),
    .D(net714),
    .RESET_B(net730),
    .Q(net805));
 sky130_fd_sc_hd__dfrtp_2 merge852 (.CLK(clknet_4_12_0_clk),
    .D(net745),
    .RESET_B(net588),
    .Q(net806));
 sky130_fd_sc_hd__dfsbp_1 merge853 (.CLK(clknet_4_15_0_clk),
    .D(net717),
    .SET_B(net616),
    .Q(net808),
    .Q_N(net807));
 sky130_fd_sc_hd__and2_0 merge854 (.A(net487),
    .B(net718),
    .X(net809));
 sky130_fd_sc_hd__dfsbp_1 merge855 (.CLK(clknet_4_11_0_clk),
    .D(net557),
    .SET_B(net675),
    .Q(net811),
    .Q_N(net810));
 sky130_fd_sc_hd__and2_0 merge856 (.A(net485),
    .B(net615),
    .X(net812));
 sky130_fd_sc_hd__dfstp_1 merge857 (.CLK(clknet_4_1_0_clk),
    .D(net749),
    .SET_B(net769),
    .Q(net964));
 sky130_fd_sc_hd__dfstp_1 merge858 (.CLK(clknet_4_15_0_clk),
    .D(net723),
    .SET_B(net493),
    .Q(net813));
 sky130_fd_sc_hd__dfstp_2 merge859 (.CLK(clknet_4_2_0_clk),
    .D(net429),
    .SET_B(net300),
    .Q(net814));
 sky130_fd_sc_hd__and2_0 merge860 (.A(net724),
    .B(net491),
    .X(net815));
 sky130_fd_sc_hd__dlrbn_1 merge861 (.D(net347),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net354),
    .Q(net817),
    .Q_N(net816));
 sky130_fd_sc_hd__dlrbn_1 merge862 (.D(net727),
    .GATE_N(clknet_4_14_0_clk),
    .RESET_B(net728),
    .Q(net819),
    .Q_N(net818));
 sky130_fd_sc_hd__dlrbp_1 merge863 (.D(net488),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net747),
    .Q(net821),
    .Q_N(net820));
 sky130_fd_sc_hd__dlrbp_1 merge864 (.D(net444),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net753),
    .Q(net823),
    .Q_N(net822));
 sky130_fd_sc_hd__dlrtn_1 merge865 (.D(net316),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net317),
    .Q(net824));
 sky130_fd_sc_hd__dlrtn_1 merge866 (.D(net674),
    .GATE_N(clknet_4_11_0_clk),
    .RESET_B(net746),
    .Q(net825));
 sky130_fd_sc_hd__dlrtn_2 merge867 (.D(net658),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net771),
    .Q(net826));
 sky130_fd_sc_hd__dlrtp_2 merge868 (.D(net620),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net710),
    .Q(net827));
 sky130_fd_sc_hd__dlrtp_1 merge869 (.D(net341),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net812),
    .Q(net828));
 sky130_fd_sc_hd__dlrtp_2 merge870 (.D(net765),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net815),
    .Q(net829));
 sky130_fd_sc_hd__edfxbp_1 merge871 (.CLK(clknet_4_4_0_clk),
    .D(net349),
    .DE(net103),
    .Q(net831),
    .Q_N(net830));
 sky130_fd_sc_hd__edfxtp_1 merge872 (.CLK(clknet_4_2_0_clk),
    .D(net318),
    .DE(net446),
    .Q(net832));
 sky130_fd_sc_hd__sdlclkp_1 merge873 (.CLK(clknet_4_6_0_clk),
    .GATE(net466),
    .SCE(net479),
    .GCLK(net833));
 sky130_fd_sc_hd__sdlclkp_2 merge874 (.CLK(clknet_4_13_0_clk),
    .GATE(net789),
    .SCE(net342),
    .GCLK(net966));
 sky130_fd_sc_hd__sdlclkp_4 merge875 (.CLK(clknet_4_14_0_clk),
    .GATE(net708),
    .SCE(net693),
    .GCLK(net834));
 sky130_fd_sc_hd__dfrbp_1 merge876 (.CLK(clknet_4_6_0_clk),
    .D(net790),
    .RESET_B(net782),
    .Q(net836),
    .Q_N(net835));
 sky130_fd_sc_hd__dfrbp_1 merge877 (.CLK(clknet_4_13_0_clk),
    .D(net741),
    .RESET_B(net809),
    .Q(net838),
    .Q_N(net837));
 sky130_fd_sc_hd__dfrtn_1 merge878 (.CLK_N(clknet_4_9_0_clk),
    .D(net564),
    .RESET_B(net561),
    .Q(net839));
 sky130_fd_sc_hd__dfrtp_2 merge879 (.CLK(clknet_4_14_0_clk),
    .D(net707),
    .RESET_B(net706),
    .Q(net840));
 sky130_fd_sc_hd__dfrtp_2 merge880 (.CLK(clknet_4_13_0_clk),
    .D(net772),
    .RESET_B(net756),
    .Q(net841));
 sky130_fd_sc_hd__dfrtp_4 merge881 (.CLK(clknet_4_1_0_clk),
    .D(net199),
    .RESET_B(net314),
    .Q(net842));
 sky130_fd_sc_hd__dfsbp_1 merge882 (.CLK(clknet_4_14_0_clk),
    .D(net571),
    .SET_B(net705),
    .Q(net844),
    .Q_N(net843));
 sky130_fd_sc_hd__dfsbp_1 merge883 (.CLK(clknet_4_6_0_clk),
    .D(net475),
    .SET_B(net495),
    .Q(net846),
    .Q_N(net845));
 sky130_fd_sc_hd__dfxbp_1 s884 (.CLK(clknet_4_4_0_clk),
    .D(net99),
    .Q(net848),
    .Q_N(net847));
 sky130_fd_sc_hd__dfxbp_2 s885 (.CLK(clknet_4_5_0_clk),
    .D(net100),
    .Q(net850),
    .Q_N(net849));
 sky130_fd_sc_hd__dfxtp_4 s886 (.CLK(clknet_4_0_0_clk),
    .D(net201),
    .Q(net851));
 sky130_fd_sc_hd__dfxtp_4 s887 (.CLK(clknet_4_1_0_clk),
    .D(net216),
    .Q(net852));
 sky130_fd_sc_hd__dfxtp_4 s888 (.CLK(clknet_4_5_0_clk),
    .D(net218),
    .Q(net853));
 sky130_fd_sc_hd__dlclkp_1 s889 (.CLK(clknet_4_5_0_clk),
    .GATE(net219),
    .GCLK(net854));
 sky130_fd_sc_hd__dlclkp_2 s890 (.CLK(clknet_4_5_0_clk),
    .GATE(net220),
    .GCLK(net855));
 sky130_fd_sc_hd__dlclkp_4 s891 (.CLK(clknet_4_5_0_clk),
    .GATE(net221),
    .GCLK(net856));
 sky130_fd_sc_hd__dlxbn_1 s892 (.D(net223),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net858),
    .Q_N(net857));
 sky130_fd_sc_hd__dlxbn_1 s893 (.D(net230),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net860),
    .Q_N(net859));
 sky130_fd_sc_hd__dlxbp_1 s894 (.D(net231),
    .GATE(clknet_4_4_0_clk),
    .Q(net862),
    .Q_N(net861));
 sky130_fd_sc_hd__dlxtn_1 s895 (.D(net233),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net863));
 sky130_fd_sc_hd__dlxtn_2 s896 (.D(net234),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net864));
 sky130_fd_sc_hd__dlxtn_1 s897 (.D(net236),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net865));
 sky130_fd_sc_hd__dlxtp_1 s898 (.D(net313),
    .GATE(clknet_4_2_0_clk),
    .Q(net866));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s899 (.D(net320),
    .SLEEP_B(clknet_4_3_0_clk),
    .Q(net867));
 sky130_fd_sc_hd__dfxbp_1 s900 (.CLK(clknet_4_7_0_clk),
    .D(net344),
    .Q(net869),
    .Q_N(net868));
 sky130_fd_sc_hd__dfxbp_1 s901 (.CLK(clknet_4_5_0_clk),
    .D(net351),
    .Q(net871),
    .Q_N(net870));
 sky130_fd_sc_hd__dfxtp_2 s902 (.CLK(clknet_4_5_0_clk),
    .D(net356),
    .Q(net965));
 sky130_fd_sc_hd__dfxtp_1 s903 (.CLK(clknet_4_7_0_clk),
    .D(net360),
    .Q(net872));
 sky130_fd_sc_hd__dfxtp_2 s904 (.CLK(clknet_4_9_0_clk),
    .D(net408),
    .Q(net873));
 sky130_fd_sc_hd__dlclkp_1 s905 (.CLK(clknet_4_9_0_clk),
    .GATE(net432),
    .GCLK(net874));
 sky130_fd_sc_hd__dlclkp_2 s906 (.CLK(clknet_4_6_0_clk),
    .GATE(net467),
    .GCLK(net875));
 sky130_fd_sc_hd__dlclkp_4 s907 (.CLK(clknet_4_3_0_clk),
    .GATE(net470),
    .GCLK(net876));
 sky130_fd_sc_hd__dlxbn_1 s908 (.D(net482),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net878),
    .Q_N(net877));
 sky130_fd_sc_hd__dlxbn_1 s909 (.D(net483),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net880),
    .Q_N(net879));
 sky130_fd_sc_hd__dlxbp_1 s910 (.D(net489),
    .GATE(clknet_4_7_0_clk),
    .Q(net882),
    .Q_N(net881));
 sky130_fd_sc_hd__dlxtn_1 s911 (.D(net490),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net883));
 sky130_fd_sc_hd__dlxtn_1 s912 (.D(net492),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net884));
 sky130_fd_sc_hd__dlxtn_4 s913 (.D(net526),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net885));
 sky130_fd_sc_hd__dlxtp_1 s914 (.D(net533),
    .GATE(clknet_4_8_0_clk),
    .Q(net886));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s915 (.D(net534),
    .SLEEP_B(clknet_4_8_0_clk),
    .Q(net887));
 sky130_fd_sc_hd__dfxbp_2 s916 (.CLK(clknet_4_9_0_clk),
    .D(net538),
    .Q(net889),
    .Q_N(net888));
 sky130_fd_sc_hd__dfxbp_2 s917 (.CLK(clknet_4_9_0_clk),
    .D(net540),
    .Q(net891),
    .Q_N(net890));
 sky130_fd_sc_hd__dfxtp_4 s918 (.CLK(clknet_4_8_0_clk),
    .D(net543),
    .Q(net892));
 sky130_fd_sc_hd__dfxtp_4 s919 (.CLK(clknet_4_9_0_clk),
    .D(net550),
    .Q(net893));
 sky130_fd_sc_hd__dfxtp_1 s920 (.CLK(clknet_4_11_0_clk),
    .D(net558),
    .Q(net894));
 sky130_fd_sc_hd__dlclkp_1 s921 (.CLK(clknet_4_11_0_clk),
    .GATE(net560),
    .GCLK(net895));
 sky130_fd_sc_hd__dlclkp_2 s922 (.CLK(clknet_4_12_0_clk),
    .GATE(net570),
    .GCLK(net896));
 sky130_fd_sc_hd__dlclkp_4 s923 (.CLK(clknet_4_12_0_clk),
    .GATE(net572),
    .GCLK(net897));
 sky130_fd_sc_hd__dlxbn_1 s924 (.D(net578),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net899),
    .Q_N(net898));
 sky130_fd_sc_hd__dlxbn_1 s925 (.D(net579),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net901),
    .Q_N(net900));
 sky130_fd_sc_hd__dlxbp_1 s926 (.D(net582),
    .GATE(clknet_4_13_0_clk),
    .Q(net903),
    .Q_N(net902));
 sky130_fd_sc_hd__dlxtn_1 s927 (.D(net584),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net904));
 sky130_fd_sc_hd__dlxtn_2 s928 (.D(net596),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net905));
 sky130_fd_sc_hd__dlxtn_1 s929 (.D(net602),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net906));
 sky130_fd_sc_hd__dlxtp_1 s930 (.D(net607),
    .GATE(clknet_4_13_0_clk),
    .Q(net907));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s931 (.D(net644),
    .SLEEP_B(clknet_4_10_0_clk),
    .Q(net908));
 sky130_fd_sc_hd__dfxbp_1 s932 (.CLK(clknet_4_10_0_clk),
    .D(net645),
    .Q(net910),
    .Q_N(net909));
 sky130_fd_sc_hd__dfxbp_1 s933 (.CLK(clknet_4_10_0_clk),
    .D(net656),
    .Q(net912),
    .Q_N(net911));
 sky130_fd_sc_hd__dfxtp_2 s934 (.CLK(clknet_4_10_0_clk),
    .D(net663),
    .Q(net913));
 sky130_fd_sc_hd__dfxtp_1 s935 (.CLK(clknet_4_11_0_clk),
    .D(net676),
    .Q(net914));
 sky130_fd_sc_hd__dfxtp_1 s936 (.CLK(clknet_4_11_0_clk),
    .D(net680),
    .Q(net915));
 sky130_fd_sc_hd__dlclkp_1 s937 (.CLK(clknet_4_11_0_clk),
    .GATE(net684),
    .GCLK(net916));
 sky130_fd_sc_hd__dlclkp_2 s938 (.CLK(clknet_4_11_0_clk),
    .GATE(net686),
    .GCLK(net917));
 sky130_fd_sc_hd__dlclkp_4 s939 (.CLK(clknet_4_11_0_clk),
    .GATE(net691),
    .GCLK(net918));
 sky130_fd_sc_hd__dlxbn_1 s940 (.D(net694),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net920),
    .Q_N(net919));
 sky130_fd_sc_hd__dlxbn_1 s941 (.D(net697),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net922),
    .Q_N(net921));
 sky130_fd_sc_hd__dlxbp_1 s942 (.D(net701),
    .GATE(clknet_4_14_0_clk),
    .Q(net924),
    .Q_N(net923));
 sky130_fd_sc_hd__dlxtn_1 s943 (.D(net702),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net925));
 sky130_fd_sc_hd__dlxtn_1 s944 (.D(net711),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net971));
 sky130_fd_sc_hd__dlxtn_1 s945 (.D(net715),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net926));
 sky130_fd_sc_hd__dlxtp_1 s946 (.D(net725),
    .GATE(clknet_4_15_0_clk),
    .Q(net927));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(in0),
    .X(net928));
 sky130_fd_sc_hd__buf_1 input2 (.A(in1),
    .X(net929));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(in10),
    .X(net930));
 sky130_fd_sc_hd__buf_1 input4 (.A(in11),
    .X(net931));
 sky130_fd_sc_hd__buf_2 input5 (.A(in12),
    .X(net932));
 sky130_fd_sc_hd__buf_4 input6 (.A(in13),
    .X(net933));
 sky130_fd_sc_hd__buf_2 input7 (.A(in14),
    .X(net934));
 sky130_fd_sc_hd__buf_6 input8 (.A(in15),
    .X(net935));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(in16),
    .X(net936));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(in17),
    .X(net937));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(in18),
    .X(net938));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(in19),
    .X(net939));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(in2),
    .X(net940));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(in20),
    .X(net941));
 sky130_fd_sc_hd__buf_2 input15 (.A(in21),
    .X(net942));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(in22),
    .X(net943));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(in23),
    .X(net944));
 sky130_fd_sc_hd__buf_2 input18 (.A(in24),
    .X(net945));
 sky130_fd_sc_hd__buf_2 input19 (.A(in3),
    .X(net946));
 sky130_fd_sc_hd__buf_12 input20 (.A(in4),
    .X(net947));
 sky130_fd_sc_hd__buf_6 input21 (.A(in5),
    .X(net948));
 sky130_fd_sc_hd__buf_2 input22 (.A(in6),
    .X(net949));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(in7),
    .X(net950));
 sky130_fd_sc_hd__buf_4 input24 (.A(in8),
    .X(net951));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(in9),
    .X(net952));
 sky130_fd_sc_hd__clkbuf_4 output26 (.A(net953),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output27 (.A(net954),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output28 (.A(net955),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output29 (.A(net996),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net957),
    .X(out13));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(clknet_1_0__leaf_net958),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output32 (.A(net1128),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output33 (.A(net960),
    .X(out16));
 sky130_fd_sc_hd__clkbuf_4 output34 (.A(net961),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output35 (.A(net962),
    .X(out19));
 sky130_fd_sc_hd__clkbuf_4 output36 (.A(net963),
    .X(out2));
 sky130_fd_sc_hd__clkbuf_4 output37 (.A(net964),
    .X(out20));
 sky130_fd_sc_hd__clkbuf_4 output38 (.A(net965),
    .X(out21));
 sky130_fd_sc_hd__clkbuf_1 output39 (.A(clknet_1_1__leaf_net966),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_1 output40 (.A(clknet_1_1__leaf_net967),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output41 (.A(net968),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output42 (.A(net1158),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output43 (.A(net970),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output44 (.A(net971),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output45 (.A(net1105),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_4 output46 (.A(net999),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_4 output47 (.A(net974),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output48 (.A(net975),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_4 fanout49 (.A(net437),
    .X(net976));
 sky130_fd_sc_hd__buf_2 fanout50 (.A(net312),
    .X(net977));
 sky130_fd_sc_hd__buf_2 fanout51 (.A(net654),
    .X(net978));
 sky130_fd_sc_hd__buf_8 fanout52 (.A(net980),
    .X(net979));
 sky130_fd_sc_hd__buf_8 fanout53 (.A(net972),
    .X(net980));
 sky130_fd_sc_hd__buf_8 fanout54 (.A(net423),
    .X(net981));
 sky130_fd_sc_hd__clkbuf_4 fanout55 (.A(net192),
    .X(net982));
 sky130_fd_sc_hd__clkbuf_4 fanout56 (.A(net187),
    .X(net983));
 sky130_fd_sc_hd__buf_8 fanout57 (.A(net385),
    .X(net984));
 sky130_fd_sc_hd__clkbuf_4 fanout58 (.A(net166),
    .X(net985));
 sky130_fd_sc_hd__buf_2 fanout59 (.A(net166),
    .X(net986));
 sky130_fd_sc_hd__clkbuf_4 fanout60 (.A(net304),
    .X(net987));
 sky130_fd_sc_hd__clkbuf_4 fanout61 (.A(net953),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_4 fanout62 (.A(net173),
    .X(net989));
 sky130_fd_sc_hd__clkbuf_4 fanout63 (.A(net279),
    .X(net990));
 sky130_fd_sc_hd__clkbuf_4 fanout64 (.A(net63),
    .X(net991));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout65 (.A(net63),
    .X(net992));
 sky130_fd_sc_hd__clkbuf_4 fanout66 (.A(net390),
    .X(net993));
 sky130_fd_sc_hd__buf_6 fanout67 (.A(net378),
    .X(net994));
 sky130_fd_sc_hd__buf_2 fanout68 (.A(net1068),
    .X(net995));
 sky130_fd_sc_hd__clkbuf_4 fanout69 (.A(net956),
    .X(net996));
 sky130_fd_sc_hd__buf_6 fanout70 (.A(net27),
    .X(net997));
 sky130_fd_sc_hd__buf_4 fanout71 (.A(net999),
    .X(net998));
 sky130_fd_sc_hd__clkbuf_4 fanout72 (.A(net973),
    .X(net999));
 sky130_fd_sc_hd__buf_4 fanout73 (.A(net139),
    .X(net1000));
 sky130_fd_sc_hd__buf_2 fanout74 (.A(net1003),
    .X(net1001));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout75 (.A(net1003),
    .X(net1002));
 sky130_fd_sc_hd__buf_2 fanout76 (.A(net1004),
    .X(net1003));
 sky130_fd_sc_hd__buf_2 fanout77 (.A(net62),
    .X(net1004));
 sky130_fd_sc_hd__buf_4 fanout78 (.A(net375),
    .X(net1005));
 sky130_fd_sc_hd__clkbuf_2 fanout79 (.A(net375),
    .X(net1006));
 sky130_fd_sc_hd__buf_4 fanout80 (.A(net25),
    .X(net1007));
 sky130_fd_sc_hd__buf_4 fanout81 (.A(net374),
    .X(net1008));
 sky130_fd_sc_hd__buf_4 fanout82 (.A(net259),
    .X(net1009));
 sky130_fd_sc_hd__clkbuf_4 fanout83 (.A(net51),
    .X(net1010));
 sky130_fd_sc_hd__buf_4 fanout84 (.A(net12),
    .X(net1011));
 sky130_fd_sc_hd__clkbuf_2 fanout85 (.A(net12),
    .X(net1012));
 sky130_fd_sc_hd__buf_8 fanout86 (.A(net1014),
    .X(net1013));
 sky130_fd_sc_hd__buf_12 fanout87 (.A(net250),
    .X(net1014));
 sky130_fd_sc_hd__clkbuf_4 fanout88 (.A(net377),
    .X(net1015));
 sky130_fd_sc_hd__clkbuf_4 fanout89 (.A(net263),
    .X(net1016));
 sky130_fd_sc_hd__buf_2 fanout90 (.A(net263),
    .X(net1017));
 sky130_fd_sc_hd__buf_4 fanout91 (.A(net133),
    .X(net1018));
 sky130_fd_sc_hd__buf_2 fanout92 (.A(net133),
    .X(net1019));
 sky130_fd_sc_hd__buf_8 fanout93 (.A(net240),
    .X(net1020));
 sky130_fd_sc_hd__buf_4 fanout94 (.A(net246),
    .X(net1021));
 sky130_fd_sc_hd__buf_6 fanout95 (.A(net2),
    .X(net1022));
 sky130_fd_sc_hd__clkbuf_4 fanout96 (.A(net387),
    .X(net1023));
 sky130_fd_sc_hd__buf_8 fanout97 (.A(net120),
    .X(net1024));
 sky130_fd_sc_hd__clkbuf_8 fanout98 (.A(net132),
    .X(net1025));
 sky130_fd_sc_hd__buf_4 fanout99 (.A(net115),
    .X(net1026));
 sky130_fd_sc_hd__clkbuf_2 max_cap100 (.A(net887),
    .X(net1027));
 sky130_fd_sc_hd__buf_4 fanout101 (.A(net886),
    .X(net1028));
 sky130_fd_sc_hd__buf_4 fanout102 (.A(net1146),
    .X(net1029));
 sky130_fd_sc_hd__clkbuf_4 fanout103 (.A(net775),
    .X(net1030));
 sky130_fd_sc_hd__buf_2 fanout104 (.A(net775),
    .X(net1031));
 sky130_fd_sc_hd__clkbuf_2 fanout105 (.A(net1033),
    .X(net1032));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout106 (.A(net1034),
    .X(net1033));
 sky130_fd_sc_hd__clkbuf_2 fanout107 (.A(net1035),
    .X(net1034));
 sky130_fd_sc_hd__clkbuf_2 fanout108 (.A(net1037),
    .X(net1035));
 sky130_fd_sc_hd__buf_4 fanout109 (.A(net1037),
    .X(net1036));
 sky130_fd_sc_hd__clkbuf_4 fanout110 (.A(net42),
    .X(net1037));
 sky130_fd_sc_hd__buf_6 fanout111 (.A(net18),
    .X(net1038));
 sky130_fd_sc_hd__clkbuf_2 fanout112 (.A(net18),
    .X(net1039));
 sky130_fd_sc_hd__buf_4 fanout113 (.A(net17),
    .X(net1040));
 sky130_fd_sc_hd__buf_4 fanout114 (.A(net4),
    .X(net1041));
 sky130_fd_sc_hd__buf_12 fanout115 (.A(net110),
    .X(net1042));
 sky130_fd_sc_hd__buf_2 fanout116 (.A(net110),
    .X(net1043));
 sky130_fd_sc_hd__buf_12 fanout117 (.A(net1045),
    .X(net1044));
 sky130_fd_sc_hd__buf_12 fanout118 (.A(net959),
    .X(net1045));
 sky130_fd_sc_hd__buf_4 fanout119 (.A(net936),
    .X(net1046));
 sky130_fd_sc_hd__buf_8 fanout120 (.A(net1048),
    .X(net1047));
 sky130_fd_sc_hd__buf_12 fanout121 (.A(net1050),
    .X(net1048));
 sky130_fd_sc_hd__buf_4 fanout122 (.A(net1050),
    .X(net1049));
 sky130_fd_sc_hd__buf_8 fanout123 (.A(net935),
    .X(net1050));
 sky130_fd_sc_hd__buf_8 fanout124 (.A(net934),
    .X(net1051));
 sky130_fd_sc_hd__clkbuf_4 fanout125 (.A(net932),
    .X(net1052));
 sky130_fd_sc_hd__buf_4 fanout126 (.A(net931),
    .X(net1053));
 sky130_fd_sc_hd__clkbuf_8 fanout127 (.A(net952),
    .X(net1054));
 sky130_fd_sc_hd__buf_4 fanout128 (.A(net950),
    .X(net1055));
 sky130_fd_sc_hd__clkbuf_4 fanout129 (.A(net950),
    .X(net1056));
 sky130_fd_sc_hd__buf_12 fanout130 (.A(net948),
    .X(net1057));
 sky130_fd_sc_hd__buf_12 fanout131 (.A(net947),
    .X(net1058));
 sky130_fd_sc_hd__buf_4 fanout132 (.A(net929),
    .X(net1059));
 sky130_fd_sc_hd__buf_4 fanout133 (.A(net946),
    .X(net1060));
 sky130_fd_sc_hd__buf_4 fanout134 (.A(net942),
    .X(net1061));
 sky130_fd_sc_hd__buf_4 fanout135 (.A(net940),
    .X(net1062));
 sky130_fd_sc_hd__buf_2 fanout136 (.A(net940),
    .X(net1063));
 sky130_fd_sc_hd__clkbuf_4 fanout137 (.A(net938),
    .X(net1064));
 sky130_fd_sc_hd__buf_8 fanout138 (.A(net937),
    .X(net1065));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net918 (.A(net918),
    .X(clknet_0_net918));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net918 (.A(clknet_0_net918),
    .X(clknet_1_0__leaf_net918));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net918 (.A(clknet_0_net918),
    .X(clknet_1_1__leaf_net918));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net917 (.A(net917),
    .X(clknet_0_net917));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net917 (.A(clknet_0_net917),
    .X(clknet_1_0__leaf_net917));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net917 (.A(clknet_0_net917),
    .X(clknet_1_1__leaf_net917));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net916 (.A(net916),
    .X(clknet_0_net916));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net916 (.A(clknet_0_net916),
    .X(clknet_1_0__leaf_net916));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net916 (.A(clknet_0_net916),
    .X(clknet_1_1__leaf_net916));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net731 (.A(net731),
    .X(clknet_0_net731));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net731 (.A(clknet_0_net731),
    .X(clknet_1_0__leaf_net731));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net731 (.A(clknet_0_net731),
    .X(clknet_1_1__leaf_net731));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net712 (.A(net712),
    .X(clknet_0_net712));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net712 (.A(clknet_0_net712),
    .X(clknet_1_0__leaf_net712));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net712 (.A(clknet_0_net712),
    .X(clknet_1_1__leaf_net712));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net720 (.A(net720),
    .X(clknet_0_net720));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net720 (.A(clknet_0_net720),
    .X(clknet_1_0__leaf_net720));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net720 (.A(clknet_0_net720),
    .X(clknet_1_1__leaf_net720));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net834 (.A(net834),
    .X(clknet_0_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net834 (.A(clknet_0_net834),
    .X(clknet_1_0__leaf_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net834 (.A(clknet_0_net834),
    .X(clknet_1_1__leaf_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net709 (.A(net709),
    .X(clknet_0_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net709 (.A(clknet_0_net709),
    .X(clknet_1_0__leaf_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net709 (.A(clknet_0_net709),
    .X(clknet_1_1__leaf_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net897 (.A(net897),
    .X(clknet_0_net897));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net897 (.A(clknet_0_net897),
    .X(clknet_1_0__leaf_net897));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net897 (.A(clknet_0_net897),
    .X(clknet_1_1__leaf_net897));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net967 (.A(net967),
    .X(clknet_0_net967));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net967 (.A(clknet_0_net967),
    .X(clknet_1_0__leaf_net967));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net967 (.A(clknet_0_net967),
    .X(clknet_1_1__leaf_net967));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net896 (.A(net896),
    .X(clknet_0_net896));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net896 (.A(clknet_0_net896),
    .X(clknet_1_0__leaf_net896));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net896 (.A(clknet_0_net896),
    .X(clknet_1_1__leaf_net896));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net895 (.A(net895),
    .X(clknet_0_net895));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net895 (.A(clknet_0_net895),
    .X(clknet_1_0__leaf_net895));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net895 (.A(clknet_0_net895),
    .X(clknet_1_1__leaf_net895));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net563 (.A(net563),
    .X(clknet_0_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net563 (.A(clknet_0_net563),
    .X(clknet_1_0__leaf_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net563 (.A(clknet_0_net563),
    .X(clknet_1_1__leaf_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net795 (.A(net795),
    .X(clknet_0_net795));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net795 (.A(clknet_0_net795),
    .X(clknet_1_0__leaf_net795));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net795 (.A(clknet_0_net795),
    .X(clknet_1_1__leaf_net795));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net562 (.A(net562),
    .X(clknet_0_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_0__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_1__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net876 (.A(net876),
    .X(clknet_0_net876));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net876 (.A(clknet_0_net876),
    .X(clknet_1_0__leaf_net876));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net876 (.A(clknet_0_net876),
    .X(clknet_1_1__leaf_net876));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net473 (.A(net473),
    .X(clknet_0_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net473 (.A(clknet_0_net473),
    .X(clknet_1_0__leaf_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net473 (.A(clknet_0_net473),
    .X(clknet_1_1__leaf_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net597 (.A(net597),
    .X(clknet_0_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net597 (.A(clknet_0_net597),
    .X(clknet_1_0__leaf_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net597 (.A(clknet_0_net597),
    .X(clknet_1_1__leaf_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net471 (.A(net471),
    .X(clknet_0_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net471 (.A(clknet_0_net471),
    .X(clknet_1_0__leaf_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net471 (.A(clknet_0_net471),
    .X(clknet_1_1__leaf_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net593 (.A(net593),
    .X(clknet_0_net593));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net593 (.A(clknet_0_net593),
    .X(clknet_1_0__leaf_net593));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net593 (.A(clknet_0_net593),
    .X(clknet_1_1__leaf_net593));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net875 (.A(net875),
    .X(clknet_0_net875));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net875 (.A(clknet_0_net875),
    .X(clknet_1_0__leaf_net875));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net875 (.A(clknet_0_net875),
    .X(clknet_1_1__leaf_net875));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net966 (.A(net966),
    .X(clknet_0_net966));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net966 (.A(clknet_0_net966),
    .X(clknet_1_0__leaf_net966));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net966 (.A(clknet_0_net966),
    .X(clknet_1_1__leaf_net966));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net721 (.A(net721),
    .X(clknet_0_net721));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net721 (.A(clknet_0_net721),
    .X(clknet_1_0__leaf_net721));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net721 (.A(clknet_0_net721),
    .X(clknet_1_1__leaf_net721));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net833 (.A(net833),
    .X(clknet_0_net833));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net833 (.A(clknet_0_net833),
    .X(clknet_1_0__leaf_net833));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net833 (.A(clknet_0_net833),
    .X(clknet_1_1__leaf_net833));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net874 (.A(net874),
    .X(clknet_0_net874));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net874 (.A(clknet_0_net874),
    .X(clknet_1_0__leaf_net874));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net874 (.A(clknet_0_net874),
    .X(clknet_1_1__leaf_net874));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net622 (.A(net622),
    .X(clknet_0_net622));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net622 (.A(clknet_0_net622),
    .X(clknet_1_0__leaf_net622));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net622 (.A(clknet_0_net622),
    .X(clknet_1_1__leaf_net622));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net856 (.A(net856),
    .X(clknet_0_net856));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net856 (.A(clknet_0_net856),
    .X(clknet_1_0__leaf_net856));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net856 (.A(clknet_0_net856),
    .X(clknet_1_1__leaf_net856));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net352 (.A(net352),
    .X(clknet_0_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net352 (.A(clknet_0_net352),
    .X(clknet_1_0__leaf_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net352 (.A(clknet_0_net352),
    .X(clknet_1_1__leaf_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net346 (.A(net346),
    .X(clknet_0_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net346 (.A(clknet_0_net346),
    .X(clknet_1_0__leaf_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net346 (.A(clknet_0_net346),
    .X(clknet_1_1__leaf_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net855 (.A(net855),
    .X(clknet_0_net855));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net855 (.A(clknet_0_net855),
    .X(clknet_1_0__leaf_net855));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net855 (.A(clknet_0_net855),
    .X(clknet_1_1__leaf_net855));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net854 (.A(net854),
    .X(clknet_0_net854));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net854 (.A(clknet_0_net854),
    .X(clknet_1_0__leaf_net854));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net854 (.A(clknet_0_net854),
    .X(clknet_1_1__leaf_net854));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net227 (.A(net227),
    .X(clknet_0_net227));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net227 (.A(clknet_0_net227),
    .X(clknet_1_0__leaf_net227));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net227 (.A(clknet_0_net227),
    .X(clknet_1_1__leaf_net227));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net958 (.A(net958),
    .X(clknet_0_net958));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net958 (.A(clknet_0_net958),
    .X(clknet_1_0__leaf_net958));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net958 (.A(clknet_0_net958),
    .X(clknet_1_1__leaf_net958));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net229 (.A(net229),
    .X(clknet_0_net229));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net229 (.A(clknet_0_net229),
    .X(clknet_1_0__leaf_net229));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net229 (.A(clknet_0_net229),
    .X(clknet_1_1__leaf_net229));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net228 (.A(net228),
    .X(clknet_0_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net228 (.A(clknet_0_net228),
    .X(clknet_1_0__leaf_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net228 (.A(clknet_0_net228),
    .X(clknet_1_1__leaf_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net222 (.A(net222),
    .X(clknet_0_net222));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net222 (.A(clknet_0_net222),
    .X(clknet_1_0__leaf_net222));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net222 (.A(clknet_0_net222),
    .X(clknet_1_1__leaf_net222));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net798 (.A(net798),
    .X(clknet_0_net798));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net798 (.A(clknet_0_net798),
    .X(clknet_1_0__leaf_net798));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net798 (.A(clknet_0_net798),
    .X(clknet_1_1__leaf_net798));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net215 (.A(net215),
    .X(clknet_0_net215));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net215 (.A(clknet_0_net215),
    .X(clknet_1_0__leaf_net215));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net215 (.A(clknet_0_net215),
    .X(clknet_1_1__leaf_net215));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net91 (.A(net91),
    .X(clknet_0_net91));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net91 (.A(clknet_0_net91),
    .X(clknet_1_0__leaf_net91));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net91 (.A(clknet_0_net91),
    .X(clknet_1_1__leaf_net91));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net97 (.A(net97),
    .X(clknet_0_net97));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net97 (.A(clknet_0_net97),
    .X(clknet_1_0__leaf_net97));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net97 (.A(clknet_0_net97),
    .X(clknet_1_1__leaf_net97));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net96 (.A(net96),
    .X(clknet_0_net96));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net96 (.A(clknet_0_net96),
    .X(clknet_1_0__leaf_net96));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net96 (.A(clknet_0_net96),
    .X(clknet_1_1__leaf_net96));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net232 (.A(net232),
    .X(clknet_0_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net232 (.A(clknet_0_net232),
    .X(clknet_1_0__leaf_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net232 (.A(clknet_0_net232),
    .X(clknet_1_1__leaf_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net95 (.A(net95),
    .X(clknet_0_net95));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net95 (.A(clknet_0_net95),
    .X(clknet_1_0__leaf_net95));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net95 (.A(clknet_0_net95),
    .X(clknet_1_1__leaf_net95));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net94 (.A(net94),
    .X(clknet_0_net94));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net94 (.A(clknet_0_net94),
    .X(clknet_1_0__leaf_net94));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net94 (.A(clknet_0_net94),
    .X(clknet_1_1__leaf_net94));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net98 (.A(net98),
    .X(clknet_0_net98));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net98 (.A(clknet_0_net98),
    .X(clknet_1_0__leaf_net98));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net98 (.A(clknet_0_net98),
    .X(clknet_1_1__leaf_net98));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net102 (.A(net102),
    .X(clknet_0_net102));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net102 (.A(clknet_0_net102),
    .X(clknet_1_0__leaf_net102));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net102 (.A(clknet_0_net102),
    .X(clknet_1_1__leaf_net102));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net797 (.A(net797),
    .X(clknet_0_net797));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net797 (.A(clknet_0_net797),
    .X(clknet_1_0__leaf_net797));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net797 (.A(clknet_0_net797),
    .X(clknet_1_1__leaf_net797));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net1156),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net1066),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net378),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net251),
    .X(net1069));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer5 (.A(net1069),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net1069),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net1069),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net111),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net1099),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net383),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net1075),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net240),
    .X(net1077));
 sky130_fd_sc_hd__clkbuf_2 rebuffer13 (.A(net423),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net1078),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net1078),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net1078),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net1194),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net21),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net1083),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net1083),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net428),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net428),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net163),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net1088),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net163),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net165),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(net165),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(net1104),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net1058),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer30 (.A(net1117),
    .X(net1095));
 sky130_fd_sc_hd__clkbuf_1 clone31 (.A(net1050),
    .X(net1096));
 sky130_fd_sc_hd__clkbuf_4 clone32 (.A(net948),
    .X(net1097));
 sky130_fd_sc_hd__clkbuf_1 clone33 (.A(net1099),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(net385),
    .X(net1099));
 sky130_fd_sc_hd__clkbuf_1 clone35 (.A(net1014),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer36 (.A(net962),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer37 (.A(net1101),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer38 (.A(net1101),
    .X(net1103));
 sky130_fd_sc_hd__clkbuf_1 clone39 (.A(net240),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer40 (.A(net980),
    .X(net1105));
 sky130_fd_sc_hd__buf_2 rebuffer41 (.A(net1105),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer42 (.A(net1106),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer43 (.A(net1106),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer44 (.A(net1112),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer45 (.A(net24),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer46 (.A(net1110),
    .X(net1111));
 sky130_fd_sc_hd__clkbuf_1 clone47 (.A(net1113),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer48 (.A(net378),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer49 (.A(net212),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer50 (.A(net1050),
    .X(net1115));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer51 (.A(net1058),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer52 (.A(net1116),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer53 (.A(net373),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer54 (.A(net507),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer55 (.A(net507),
    .X(net1120));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer56 (.A(net507),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer57 (.A(net1121),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer58 (.A(net400),
    .X(net1123));
 sky130_fd_sc_hd__clkbuf_1 rebuffer59 (.A(net400),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer60 (.A(net1124),
    .X(net1125));
 sky130_fd_sc_hd__clkbuf_4 clone61 (.A(net1045),
    .X(net1126));
 sky130_fd_sc_hd__clkbuf_1 clone62 (.A(net1048),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer63 (.A(net1045),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer64 (.A(net569),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer65 (.A(net569),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer66 (.A(net984),
    .X(net1131));
 sky130_fd_sc_hd__clkbuf_1 clone67 (.A(net980),
    .X(net1132));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer68 (.A(net654),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer69 (.A(net1133),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer70 (.A(net1134),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net851),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net781),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net886),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net762),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net927),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net893),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net907),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net964),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net637),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net926),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net866),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net842),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net909),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net910),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net791),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net828),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net908),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net911),
    .X(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A0 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_D1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_S1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_B (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c30_A (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A2 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c25_X (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c49_A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_C (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_A (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_A1 (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c35_X (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A0 (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_C1 (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_B (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_Q (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A0 (.DIODE(net1184));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A1 (.DIODE(net1183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_D1 (.DIODE(net1191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A3 (.DIODE(net1191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_B (.DIODE(net1191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A (.DIODE(net1191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B (.DIODE(net1191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A (.DIODE(net1191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net1191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A3 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_C1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_X (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_B (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_B1 (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_X (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c49_C1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_X (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A0 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_X (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer8_A (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_SCE (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_C (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_B (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_X (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c659_A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A0 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A3 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_C1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_S1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_X (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_X (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer17_A (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A1 (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_B (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_S1 (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_X (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A3 (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_C1 (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_B (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A3 (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A1 (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_B (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_B (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_X (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_C1 (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A1 (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_B (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_B (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_X (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A1 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_A1 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_SCD (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A3 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_B (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A2 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A0 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_X (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_B (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_B (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_S1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_X (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout97_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A0 (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A3 (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_X (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_D1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_C (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_X (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_D1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_C_N (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_X (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_A3 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_D1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A0 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_C (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_C1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_X (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c55_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c39_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_X (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_A3 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_X (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_X (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_D1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_C_N (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_C (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_X (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A3 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_D1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_X (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A0 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_C (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A3 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_X (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_C (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_D_N (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_D1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_X (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_A0 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c39_X (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A0 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_B (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_X (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c649_A0 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A0 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A3 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_D1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_X (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A0 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A0 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A0 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S0 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_X (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S0 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A0 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_D1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_C_N (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_X (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_D_N (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_D1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_C_N (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_X (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A0 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A3 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_X (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A0 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_SCD (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_C1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_X (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A0 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_X (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A0 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_S0 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_X (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_D_N (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_D_N (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_X (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_X (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A0 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_C1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_D1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_X (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S0 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A3 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A3 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_C_N (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_X (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A0 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A3 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_D1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_X (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_B (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A0 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_X (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_C (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S0 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_X (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A0 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_S1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S0 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_X (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c658_A0 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_A3 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_X (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A3 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A0 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A3 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_X (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A0 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A0 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A3 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A3 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A3 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_C1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_X (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_A0 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_X (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_X (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A3 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_D1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_X (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_X (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_C1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A3 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_SCD (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A3 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_C_N (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_X (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A0 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_X (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A0 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_C1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_C1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_X (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_S0 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A0 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S0 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_C1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_C (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_C (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_X (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_X (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_X (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout56_A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_S0 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_X (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A3 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A3 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_C1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_C1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_Q_N (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_C (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c44_X (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_C1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c658_S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c652_A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_Q (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout55_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_A0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_X (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_Q (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A0 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_S0 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_X (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_C1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A3 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c27_X (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c45_X (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_C (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A0 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S0 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_D1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_SCD (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_C1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_C1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_S0 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_X (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c49_D1 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer18_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_B (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c46_X (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A0 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A3 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_C1 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c47_X (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_D1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_C (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c657_A0 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_X (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_S1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_B (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_C1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S0 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A0 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c52_B1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c48_X (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_C (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_X (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone39_A (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer12_A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout93_A (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A3 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A0 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_C_N (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_X (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A0 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S0 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_S1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_X (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A0 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S0 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_C_N (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_X (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A0 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_X (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout94_A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c643_A3 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_C1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_X (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_X (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_C_N (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_X (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c50_X (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer4_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_C_N (.DIODE(net1185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A3 (.DIODE(net1185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_C1 (.DIODE(net1185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_B1 (.DIODE(net1185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A0 (.DIODE(net1185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_X (.DIODE(net1185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_S0 (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A3 (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_D1 (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A1 (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A3 (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A0 (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A1 (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_X (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_C1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_A (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_C_N (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A1 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_X (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S0 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A0 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A0 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S0 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_X (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S0 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A1 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A2 (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A2 (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A3 (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A2 (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_X (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_X (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c653_A3 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c648_A0 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A0 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_S1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_S1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_C (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_X (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_C (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_X (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A3 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A0 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_X (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_D1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_X (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A0 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c52_X (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A0 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_S0 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_X (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_SCD (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_C1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_C1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_X (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A0 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_C1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_B1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_X (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A0 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S0 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_X (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_S0 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_C1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_X (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A3 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c53_X (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c45_A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_D_N (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_D1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A2 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A0 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_S0 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_B (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_X (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A2 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_B1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A2 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A0 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_C (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_X (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A0 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A2 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S0 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_X (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A2 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_C (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_X (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_B1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A0 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A3 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A3 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A3 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_X (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_A0 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A3 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_C (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_X (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_C1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A0 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_X (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A0 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c56_B (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c54_X (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c45_A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_RESET_B (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A0 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_S1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A0 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_X (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A0 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_X (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_A0 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_S0 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_X (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A0 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A3 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_X (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c53_B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_A3 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c30_B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c28_X (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_X (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c57_X (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c50_C1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A3 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A0 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_C_N (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_A2 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_S0 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A2 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A2 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_X (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A3 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A0 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S0 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A3 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A2 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_B1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A3 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_X (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_A3 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A3 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_B1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A0 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_B1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_X (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_A0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_X (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_A0 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_S0 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_X (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_C_N (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A3 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c58_X (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c52_A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c60_X (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S0 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c48_B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A3 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c61_X (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c46_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_C (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A2 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_C1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_S0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A3 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A2 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_X (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A0 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A3 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_X (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A0 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_C_N (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_X (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S1 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_X (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_A (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_A (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_X (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A0 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_X (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_X (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c51_B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c50_B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c48_C_N (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c47_B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A3 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A0 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A0 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S0 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A3 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A0 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_X (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A0 (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A1 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_X (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_SCD (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_B (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_B (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A1 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_X (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A0 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S0 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_C (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_X (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A1 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_X (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_X (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_RESET_B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c47_A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_X (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_X (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_C1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_B (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_X (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A3 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A2 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A0 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A0 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_C (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_X (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_D1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_X (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A0 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A3 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A3 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_X (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_S1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_X (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A0 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_B1 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_B (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_D1 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_X (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A1 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A1 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A1 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_X (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A3 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_X (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_S0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_X (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_S1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A2 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_X (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_A2 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_A0 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A3 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A3 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_X (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_X (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_C1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A3 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_C_N (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_Q_N (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_RESET_B (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_Q (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A3 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_X (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_A3 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_A1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_B (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_C_N (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_X (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_X (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A1 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_X (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout49_A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A0 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_A0 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_X (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A0 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_C_N (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A0 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_X (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A0 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S0 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A2 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A2 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_SET_B (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_X (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S0 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_X (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_X (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A3 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge850_RESET_B (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_X (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_c643_A0 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S0 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_X (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_A0 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S0 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A3 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S0 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_X (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_c650_A0 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A3 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_A2 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_A3 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A2 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_X (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_A0 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_S1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_X (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_B (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_X (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S0 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_C_N (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_X (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A3 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_X (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A0 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_SET_B (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_X (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_C (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_X (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A3 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A0 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A3 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_C (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A1 (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A0 (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_X (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A2 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S0 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A2 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A2 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_B (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_X (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A3 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A0 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S0 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A0 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A1 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A3 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_B (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_C (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_X (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_C1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_X (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S0 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A3 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A3 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A0 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_SCE (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_X (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A0 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A3 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S1 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A2 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S0 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A3 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_S0 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S1 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_Q_N (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_A1 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_S0 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_A2 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A1 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S0 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S1 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A2 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_Q (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_B1 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A1 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A3 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_S1 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A0 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_X (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_S0 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A1 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A0 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A1 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A3 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A1 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_X (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_D1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_S0 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_S0 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_S0 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_Q_N (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A0 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A1 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A3 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A2 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A1 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_X (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A0 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A0 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A2 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_X (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_B (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_X (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A0 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_S0 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c650_A1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S0 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A2 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S0 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_S0 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_X (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A2 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A1 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A0 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A3 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A3 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_X (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_X (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A3 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_S1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_X (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A0 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A0 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S0 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A3 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_X (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A3 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S0 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A3 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S0 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_X (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_B (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_X (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A0 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c659_A0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_X (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A3 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A1 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A3 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_X (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer65_A (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer64_A (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A0 (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_X (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A0 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_X (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_A2 (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c652_S0 (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A3 (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_S0 (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A3 (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_B1 (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_B1 (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A0 (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_X (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_S0 (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A0 (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A3 (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_A1 (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_C_N (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A0 (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_A (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A0 (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A2 (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c35_C_N (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A1 (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c31_X (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_B1 (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_D1 (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_S0 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_X (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_D (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_X (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A2 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A1 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A3 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_S0 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_X (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A0 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A2 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A3 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A1 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_X (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A3 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A3 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A2 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A2 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_Q_N (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A0 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A1 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A2 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_B (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_Q (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_X (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_S0 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_S0 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A3 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_X (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_X (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A0 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_S1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A0 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A3 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A3 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A0 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_X (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A0 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_X (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A0 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_X (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_X (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A2 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S0 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A3 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_X (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_X (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_X (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c35_B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c57_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_C (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c32_X (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_D1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_X (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A3 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_X (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_Q (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_D (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_X (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_Q_N (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_X (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold85_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_Q (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S0 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_D_N (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_C_N (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_D1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_Q (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A3 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S0 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S0 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S0 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A2 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge848_Q (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_S0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A3 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge850_Q (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_S0 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_C1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A3 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_A3 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_X (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_Q (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S0 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_A2 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_Q (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S0 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_D1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_C (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_D_N (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_Q (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A3 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A3 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S1 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_D1 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_C1 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_Q (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A3 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A3 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_Q (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A2 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A3 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_S1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_Q (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A2 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A2 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c657_A3 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_S0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_Q (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_A3 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_Q (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_A3 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_A3 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_Q (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_D1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_B1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_Q (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S0 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_S1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S0 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S0 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_A0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_S0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_S1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold82_A (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_Q (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_D1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_C1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_S0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_D1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_S1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_Q (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_S1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_Q_N (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_S1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_S0 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_SET_B (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A3 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_D1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_X (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_Q (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c648_A3 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_A3 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_S0 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_S1 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold71_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_Q (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S0 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_D1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_D1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_D1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_Q (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_S0 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_S0 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A3 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_S1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_S1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_S0 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_Q (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_A3 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_S1 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A2 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_S1 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_S0 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_S1 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_S1 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_S0 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_S1 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_S1 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_S0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_D1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_C (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_X (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_Q (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c653_S1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_S1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_Q (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_S0 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_S0 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_Q (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_A3 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_S0 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_S1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_Q (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_S0 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_S1 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_S0 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_S1 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_S1 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S0 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_S1 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold81_A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_S1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_Q (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_Q (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A3 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_D1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_Q (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_S0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c645_S0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c643_S1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_Q (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S0 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_S0 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_S1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_S1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_S1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_Q_N (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S0 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_Q (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_S0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_S1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A3 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_SCE (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_C_N (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_X (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_Q (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_S1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_Q (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_S0 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold76_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_Q (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_Q (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_S0 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c48_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c39_B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_X (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_Q (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S0 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold87_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_Q (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_S0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_S1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_Q (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_S1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S0 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A3 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_S0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_X (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c50_A1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c45_C1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_B (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A3 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c55_A (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S0 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_B1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A0 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_C1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A2 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A0 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_B (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_B (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_B (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_B1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_B (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A0 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c61_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_B (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c46_A2 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_B1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_C1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_B (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c58_B (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c25_B (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S0 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_C1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A0 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_B (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_S0 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_A1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_B1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_B (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_S0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_A (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_C1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c25_A (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_B (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_B (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_A3 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_B (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A2 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_B (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A2 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c27_A (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A2 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A0 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S0 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c643_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone32_A (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A2 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_B (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_B (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A3 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_C (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c57_B (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_S0 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_D_N (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_B1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_B (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_output26_A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_X (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_output27_A (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_B (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_SCD (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_X (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_output28_A (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_Q (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout69_A (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_X (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c652_A3 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_output33_A (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_RESET_B (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_X (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer36_A (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_A (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_D_N (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_C_N (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_X (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_output36_A (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_C1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A2 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_X (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold78_A (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_output37_A (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_Q (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A3 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S0 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_output38_A (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_Q (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_S1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c650_S1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_S0 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_S1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_S1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_S1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_S1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_output41_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_Q (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_output42_A (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_X (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A1 (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A1 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A1 (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_D_N (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA_output43_A (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_S0 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A0 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_C_N (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_S0 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_C1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_C (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_C1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_output48_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_Q (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_S0 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_S0 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_S1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout49_X (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_A2 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A3 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_SET_B (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A3 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_D1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_C1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A2 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_C1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_B1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_X (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A2 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A2 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A2 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A3 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A0 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_B1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A2 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A2 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A3 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_X (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S0 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A3 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S0 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A3 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_S1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A2 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A3 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_X (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A3 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A3 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A3 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_S1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S0 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_SCD (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A3 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout55_X (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c653_A2 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_D1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A0 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A2 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A2 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_S0 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout56_X (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A0 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A3 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_S0 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A3 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A3 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_B1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_D (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_S1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_X (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A2 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A2 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_D1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_B1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_D1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_C1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_C1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A2 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_B1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_X (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S0 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S0 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A3 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S0 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_X (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A2 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A0 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_S0 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A2 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A2 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_C1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_C1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A2 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_X (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_A2 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A3 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A2 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A2 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_X (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A3 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A2 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A2 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_C_N (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A2 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_C1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A3 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A2 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_X (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A3 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_B1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A3 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_B1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A3 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_C (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A2 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A2 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_X (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_B1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_B1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_A3 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_C (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_B1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_B1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_C1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_D1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_C1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_B1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_X (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A0 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_B1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_X (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_A3 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c649_A3 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A3 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_B (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout69_X (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_output29_A (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_B (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_C (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_D1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_B1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_A3 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_D1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_X (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_S0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_D1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_SCE (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_S1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_C1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_C (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A3 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_X (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A3 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A0 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_S1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_B (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_D1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_D1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_C1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_D_N (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_X (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_output46_A (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_A (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_X (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_C1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_S0 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_C1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_X (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_B1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_S1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_A (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_D1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_A (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_A (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_X (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c650_A3 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c648_A1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_S0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_C1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_X (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_S1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_C_N (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A0 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A3 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A3 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_S0 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A3 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_C (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_X (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S0 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S0 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c52_C1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c44_A (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A2 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_S1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_D1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_X (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A3 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_S0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_B (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A3 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_X (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A2 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A2 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_S0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_S0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_C (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A2 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_C (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A2 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_X (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_S0 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_S0 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_S1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_A1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A0 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_S0 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_X (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S0 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_C (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_C (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_A1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_C1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_C1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S0 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_S0 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_X (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A2 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S0 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A2 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S0 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone35_A (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_X (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c658_A2 (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A0 (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A1 (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S0 (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_A (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_X (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S0 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S0 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_C_N (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_D1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A3 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_X (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_C1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_B1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_D1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_C1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_S0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A3 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A3 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A3 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_X (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_S1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A3 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A3 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_X (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_B (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_S1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_X (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A0 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout94_X (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_S0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A2 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_SET_B (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_C (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_X (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_C (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_B1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_C (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_A (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c61_C (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c32_A (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A2 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_B (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c31_B (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_C (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_X (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_C_N (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_D1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A3 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout97_X (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_C1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_C1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_B1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_B1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A2 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_B1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_A1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_X (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_D1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_A0 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_C1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_S0 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_C (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_C (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_D_N (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_X (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A3 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_C (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S0 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_C (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_B (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A3 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_D1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_B (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap100_X (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S0 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S0 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_X (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_S1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_S1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_S1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_S0 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_S0 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_S0 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_S1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout102_X (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_S1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S0 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_D1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_S1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_S1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_S1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_X (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_D_N (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A3 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_D1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_D1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_D_N (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_D1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_D1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_SET_B (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_D1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_X (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A3 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_D1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_S1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_X (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_S1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_D1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A2 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_D_N (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_X (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A3 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_A1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_S0 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S0 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S0 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_D1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_D1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_D_N (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_X (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_S0 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_S1 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_S0 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_X (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c54_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_A2 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_D1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_S0 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c33_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_S0 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_X (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A2 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S0 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A1 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A3 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_X (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_S0 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_A2 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_D1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S0 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_B1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_C1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_S0 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A2 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_X (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c47_C1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A3 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_D1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_D_N (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_D1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_C_N (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_A0 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_X (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A2 (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A2 (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_C_N (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_D1 (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_S0 (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_C1 (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_X (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_D1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_B1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_X (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_D1 (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer63_A (.DIODE(net1198));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone61_A (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_X (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_S1 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_C1 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A3 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A3 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_C (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_X (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A1 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A3 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A1 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_S1 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A3 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c50_D1 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_B (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_X (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_S1 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c55_C (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c46_S1 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c35_D_N (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone62_A (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_X (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_A (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_D1 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_C (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_D1 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_C1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_X (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A0 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_A1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A2 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_B1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_D1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A3 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S0 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_S0 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer50_A (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone31_A (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_X (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_A0 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c657_A1 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_X (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A3 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A0 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c51_A (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_C1 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A1 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S1 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_X (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A1 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A3 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A1 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A1 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_D (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A0 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_A (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_C1 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S0 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_X (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c645_A0 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S0 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_A1 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A1 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A3 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S0 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A2 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A1 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_D1 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_X (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S1 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_D_N (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c643_A1 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A1 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_A3 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S0 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A1 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_X (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A3 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_S1 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_S1 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A3 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_C (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c33_A (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_C_N (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_S0 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_D1 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_X (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S0 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A1 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A1 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A3 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S0 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A0 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_X (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A3 (.DIODE(net1193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A (.DIODE(net1193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A (.DIODE(net1193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A3 (.DIODE(net1193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A (.DIODE(net1193));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer51_A (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer29_A (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_X (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A0 (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_A (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_B (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_S1 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A3 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A3 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A0 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_A (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_S0 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c28_A (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_B (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_X (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A1 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A3 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A3 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A1 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_C (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_B1 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A1 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_C (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_X (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_A1 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_A1 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c56_A (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A3 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S1 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A3 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_S0 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A1 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_X (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A3 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_A (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c52_D1 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_C (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_C (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_A (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_S1 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_C1 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_X (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A1 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_S0 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_A3 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_X (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A2 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_B (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_SCE (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_C (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_A (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c54_A (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c50_A2 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c49_A1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_S0 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_X (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_S1 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A3 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A0 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_C_N (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A3 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_A (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S0 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_B (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge847_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge864_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_SLEEP_B (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge828_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s908_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s905_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge848_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_SLEEP_B (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s933_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_S1 (.DIODE(clknet_1_0__leaf_net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c645_S1 (.DIODE(clknet_1_0__leaf_net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net896_X (.DIODE(clknet_1_0__leaf_net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(clknet_1_1__leaf_net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_output39_A (.DIODE(clknet_1_1__leaf_net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net966_X (.DIODE(clknet_1_1__leaf_net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A1 (.DIODE(clknet_1_1__leaf_net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c649_A2 (.DIODE(clknet_1_1__leaf_net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net227_X (.DIODE(clknet_1_1__leaf_net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_S1 (.DIODE(clknet_1_0__leaf_net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A (.DIODE(clknet_1_0__leaf_net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net798_X (.DIODE(clknet_1_0__leaf_net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_A (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer3_X (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_A (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_A2 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer6_A (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer5_A (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_S1 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer4_X (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_A0 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A0 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A2 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer8_X (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer16_A (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer15_A (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A2 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer14_A (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer13_X (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer24_A (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer23_X (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_A1 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer24_X (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A0 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer25_X (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer27_X (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_SCE (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S0 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_C1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_C1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_A2 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone31_X (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A0 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_A3 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A0 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S1 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A2 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone32_X (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A3 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A3 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A3 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A2 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A1 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone33_X (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A0 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_S1 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_C (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A3 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_B (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone35_X (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer38_A (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer37_A (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer36_X (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer28_A (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A2 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_B (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S1 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone39_X (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer41_A (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_A (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer40_X (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer43_A (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer42_A (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer41_X (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_C1 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A3 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_D1 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_S0 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone61_X (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c48_D_N (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_B (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_C1 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_C (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S1 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone62_X (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A3 (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A2 (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_S0 (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_S0 (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A2 (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone67_X (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout102_A (.DIODE(net1146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A3 (.DIODE(net1146));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold81_X (.DIODE(net1146));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net718));
 sky130_fd_sc_hd__mux4_1 clone1 (.A0(net44),
    .A1(net1011),
    .A2(net53),
    .A3(net1060),
    .S0(net46),
    .S1(net55),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer31 (.A(net255),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(net1155),
    .X(net1156));
 sky130_fd_sc_hd__mux4_1 clone34 (.A0(net1),
    .A1(net36),
    .A2(net939),
    .A3(net15),
    .S0(net31),
    .S1(net1047),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer35 (.A(net969),
    .X(net1158));
 sky130_fd_sc_hd__buf_2 rebuffer39 (.A(net1158),
    .X(net1159));
 sky130_fd_sc_hd__and2_1 clone40 (.A(net1194),
    .B(net116),
    .X(net1160));
 sky130_fd_sc_hd__or4bb_1 clone41 (.A(net1021),
    .B(net252),
    .C_N(net962),
    .D_N(net1013),
    .X(net1161));
 sky130_fd_sc_hd__or4bb_1 clone42 (.A(net5),
    .B(net7),
    .C_N(net1047),
    .D_N(net6),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer47 (.A(net258),
    .X(net1163));
 sky130_fd_sc_hd__or4bb_1 clone48 (.A(net256),
    .B(net1104),
    .C_N(net242),
    .D_N(net951),
    .X(net1164));
 sky130_fd_sc_hd__and2_1 clone49 (.A(net5),
    .B(net1022),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer61 (.A(net382),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer62 (.A(net1166),
    .X(net1167));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer67 (.A(net384),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer71 (.A(net1168),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer72 (.A(net1169),
    .X(net1170));
 sky130_fd_sc_hd__and3_1 clone73 (.A(net1042),
    .B(net1054),
    .C(net1060),
    .X(net1171));
 sky130_fd_sc_hd__and2_1 clone74 (.A(net123),
    .B(net1197),
    .X(net1172));
 sky130_fd_sc_hd__mux4_1 clone75 (.A0(net307),
    .A1(net567),
    .A2(net1009),
    .A3(net1194),
    .S0(net811),
    .S1(net893),
    .X(net1173));
 sky130_fd_sc_hd__and2_1 clone76 (.A(net109),
    .B(net107),
    .X(net1174));
 sky130_fd_sc_hd__and2_1 clone77 (.A(net116),
    .B(net108),
    .X(net1175));
 sky130_fd_sc_hd__and2_1 clone78 (.A(net111),
    .B(net1042),
    .X(net1176));
 sky130_fd_sc_hd__and2_1 clone79 (.A(net115),
    .B(net1043),
    .X(net1177));
 sky130_fd_sc_hd__and2_1 clone80 (.A(net1183),
    .B(net1044),
    .X(net1178));
 sky130_fd_sc_hd__and2_1 clone81 (.A(net1044),
    .B(net939),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer82 (.A(net58),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer83 (.A(net1180),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer84 (.A(net1180),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer85 (.A(net106),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer86 (.A(net1183),
    .X(net1184));
 sky130_fd_sc_hd__a2111o_1 clone87 (.A1(net113),
    .A2(net245),
    .B1(net249),
    .C1(net1013),
    .D1(net1126),
    .X(net1185));
 sky130_fd_sc_hd__clkbuf_1 clone88 (.A(net947),
    .X(net1186));
 sky130_fd_sc_hd__clkbuf_1 clone89 (.A(net110),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer90 (.A(net57),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer91 (.A(net1188),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer92 (.A(net1189),
    .X(net1190));
 sky130_fd_sc_hd__and3_1 clone93 (.A(net1047),
    .B(net1051),
    .C(net951),
    .X(net1191));
 sky130_fd_sc_hd__clkbuf_1 clone94 (.A(net959),
    .X(net1192));
 sky130_fd_sc_hd__clkbuf_1 clone95 (.A(net948),
    .X(net1193));
 sky130_fd_sc_hd__and2_1 clone96 (.A(net109),
    .B(net107),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer97 (.A(net109),
    .X(net1195));
 sky130_fd_sc_hd__clkbuf_1 clone98 (.A(net250),
    .X(net1196));
 sky130_fd_sc_hd__clkbuf_1 clone99 (.A(net1198),
    .X(net1197));
 sky130_fd_sc_hd__clkbuf_1 clone100 (.A(net959),
    .X(net1198));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
