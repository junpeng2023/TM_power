module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in62,
    in63,
    in64,
    in65,
    in66,
    in67,
    in68,
    in69,
    in7,
    in70,
    in71,
    in72,
    in73,
    in74,
    in75,
    in76,
    in77,
    in78,
    in79,
    in8,
    in80,
    in81,
    in82,
    in83,
    in84,
    in85,
    in86,
    in87,
    in88,
    in89,
    in9,
    in90,
    in91,
    in92,
    in93,
    in94,
    in95,
    in96,
    in97,
    in98,
    in99,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out62,
    out63,
    out64,
    out65,
    out66,
    out67,
    out68,
    out69,
    out7,
    out70,
    out71,
    out72,
    out73,
    out74,
    out75,
    out76,
    out77,
    out78,
    out79,
    out8,
    out80,
    out81,
    out82,
    out83,
    out84,
    out85,
    out86,
    out87,
    out88,
    out89,
    out9,
    out90,
    out91,
    out92,
    out93,
    out94,
    out95,
    out96,
    out97,
    out98,
    out99,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in62;
 input in63;
 input in64;
 input in65;
 input in66;
 input in67;
 input in68;
 input in69;
 input in7;
 input in70;
 input in71;
 input in72;
 input in73;
 input in74;
 input in75;
 input in76;
 input in77;
 input in78;
 input in79;
 input in8;
 input in80;
 input in81;
 input in82;
 input in83;
 input in84;
 input in85;
 input in86;
 input in87;
 input in88;
 input in89;
 input in9;
 input in90;
 input in91;
 input in92;
 input in93;
 input in94;
 input in95;
 input in96;
 input in97;
 input in98;
 input in99;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out62;
 output out63;
 output out64;
 output out65;
 output out66;
 output out67;
 output out68;
 output out69;
 output out7;
 output out70;
 output out71;
 output out72;
 output out73;
 output out74;
 output out75;
 output out76;
 output out77;
 output out78;
 output out79;
 output out8;
 output out80;
 output out81;
 output out82;
 output out83;
 output out84;
 output out85;
 output out86;
 output out87;
 output out88;
 output out89;
 output out9;
 output out90;
 output out91;
 output out92;
 output out93;
 output out94;
 output out95;
 output out96;
 output out97;
 output out98;
 output out99;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net764;
 wire clknet_1_0__leaf_net764;
 wire clknet_1_1__leaf_net764;
 wire clknet_0_net650;
 wire clknet_1_0__leaf_net650;
 wire clknet_1_1__leaf_net650;
 wire clknet_0_net526;
 wire clknet_1_0__leaf_net526;
 wire clknet_1_1__leaf_net526;
 wire clknet_0_net527;
 wire clknet_1_0__leaf_net527;
 wire clknet_1_1__leaf_net527;
 wire clknet_0_net525;
 wire clknet_1_0__leaf_net525;
 wire clknet_1_1__leaf_net525;
 wire clknet_0_net547;
 wire clknet_1_0__leaf_net547;
 wire clknet_1_1__leaf_net547;
 wire clknet_0_net879;
 wire clknet_1_0__leaf_net879;
 wire clknet_1_1__leaf_net879;
 wire clknet_0_net436;
 wire clknet_1_0__leaf_net436;
 wire clknet_1_1__leaf_net436;
 wire clknet_0_net891;
 wire clknet_1_0__leaf_net891;
 wire clknet_1_1__leaf_net891;
 wire clknet_0_net423;
 wire clknet_1_0__leaf_net423;
 wire clknet_1_1__leaf_net423;
 wire clknet_0_net427;
 wire clknet_1_0__leaf_net427;
 wire clknet_1_1__leaf_net427;
 wire clknet_0_net878;
 wire clknet_1_0__leaf_net878;
 wire clknet_1_1__leaf_net878;
 wire clknet_0_net422;
 wire clknet_1_0__leaf_net422;
 wire clknet_1_1__leaf_net422;
 wire clknet_0_net424;
 wire clknet_1_0__leaf_net424;
 wire clknet_1_1__leaf_net424;
 wire clknet_0_net746;
 wire clknet_1_0__leaf_net746;
 wire clknet_1_1__leaf_net746;
 wire clknet_0_net416;
 wire clknet_1_0__leaf_net416;
 wire clknet_1_1__leaf_net416;
 wire clknet_0_net728;
 wire clknet_1_0__leaf_net728;
 wire clknet_1_1__leaf_net728;
 wire clknet_0_net887;
 wire clknet_1_0__leaf_net887;
 wire clknet_1_1__leaf_net887;
 wire clknet_0_net365;
 wire clknet_1_0__leaf_net365;
 wire clknet_1_1__leaf_net365;
 wire clknet_0_net496;
 wire clknet_1_0__leaf_net496;
 wire clknet_1_1__leaf_net496;
 wire clknet_0_net727;
 wire clknet_1_0__leaf_net727;
 wire clknet_1_1__leaf_net727;
 wire clknet_0_net466;
 wire clknet_1_0__leaf_net466;
 wire clknet_1_1__leaf_net466;
 wire clknet_0_net484;
 wire clknet_1_0__leaf_net484;
 wire clknet_1_1__leaf_net484;
 wire clknet_0_net368;
 wire clknet_1_0__leaf_net368;
 wire clknet_1_1__leaf_net368;
 wire clknet_0_net376;
 wire clknet_1_0__leaf_net376;
 wire clknet_1_1__leaf_net376;
 wire clknet_0_net364;
 wire clknet_1_0__leaf_net364;
 wire clknet_1_1__leaf_net364;
 wire clknet_0_net382;
 wire clknet_1_0__leaf_net382;
 wire clknet_1_1__leaf_net382;
 wire clknet_0_net398;
 wire clknet_1_0__leaf_net398;
 wire clknet_1_1__leaf_net398;
 wire clknet_0_net384;
 wire clknet_1_0__leaf_net384;
 wire clknet_1_1__leaf_net384;
 wire clknet_0_net363;
 wire clknet_1_0__leaf_net363;
 wire clknet_1_1__leaf_net363;
 wire clknet_0_net361;
 wire clknet_1_0__leaf_net361;
 wire clknet_1_1__leaf_net361;
 wire clknet_0_net726;
 wire clknet_1_0__leaf_net726;
 wire clknet_1_1__leaf_net726;
 wire clknet_0_net396;
 wire clknet_1_0__leaf_net396;
 wire clknet_1_1__leaf_net396;
 wire clknet_0_net506;
 wire clknet_1_0__leaf_net506;
 wire clknet_1_1__leaf_net506;
 wire clknet_0_net532;
 wire clknet_1_0__leaf_net532;
 wire clknet_1_1__leaf_net532;
 wire clknet_0_net499;
 wire clknet_1_0__leaf_net499;
 wire clknet_1_1__leaf_net499;
 wire clknet_0_net875;
 wire clknet_1_0__leaf_net875;
 wire clknet_1_1__leaf_net875;
 wire clknet_0_net383;
 wire clknet_1_0__leaf_net383;
 wire clknet_1_1__leaf_net383;
 wire clknet_0_net278;
 wire clknet_1_0__leaf_net278;
 wire clknet_1_1__leaf_net278;
 wire clknet_0_net300;
 wire clknet_1_0__leaf_net300;
 wire clknet_1_1__leaf_net300;
 wire clknet_0_net293;
 wire clknet_1_0__leaf_net293;
 wire clknet_1_1__leaf_net293;
 wire clknet_0_net314;
 wire clknet_1_0__leaf_net314;
 wire clknet_1_1__leaf_net314;
 wire clknet_0_net316;
 wire clknet_1_0__leaf_net316;
 wire clknet_1_1__leaf_net316;
 wire clknet_0_net303;
 wire clknet_1_0__leaf_net303;
 wire clknet_1_1__leaf_net303;
 wire clknet_0_net912;
 wire clknet_1_0__leaf_net912;
 wire clknet_1_1__leaf_net912;
 wire clknet_0_net277;
 wire clknet_1_0__leaf_net277;
 wire clknet_1_1__leaf_net277;
 wire clknet_0_net709;
 wire clknet_1_0__leaf_net709;
 wire clknet_1_1__leaf_net709;
 wire clknet_0_net489;
 wire clknet_1_0__leaf_net489;
 wire clknet_1_1__leaf_net489;
 wire clknet_0_net478;
 wire clknet_1_0__leaf_net478;
 wire clknet_1_1__leaf_net478;
 wire clknet_0_net275;
 wire clknet_1_0__leaf_net275;
 wire clknet_1_1__leaf_net275;
 wire clknet_0_net708;
 wire clknet_1_0__leaf_net708;
 wire clknet_1_1__leaf_net708;
 wire clknet_0_net335;
 wire clknet_1_0__leaf_net335;
 wire clknet_1_1__leaf_net335;
 wire clknet_0_net907;
 wire clknet_1_0__leaf_net907;
 wire clknet_1_1__leaf_net907;
 wire clknet_0_net894;
 wire clknet_1_0__leaf_net894;
 wire clknet_1_1__leaf_net894;
 wire clknet_0_net330;
 wire clknet_1_0__leaf_net330;
 wire clknet_1_1__leaf_net330;
 wire clknet_0_net339;
 wire clknet_1_0__leaf_net339;
 wire clknet_1_1__leaf_net339;
 wire clknet_0_net338;
 wire clknet_1_0__leaf_net338;
 wire clknet_1_1__leaf_net338;
 wire clknet_0_net262;
 wire clknet_1_0__leaf_net262;
 wire clknet_1_1__leaf_net262;
 wire clknet_0_net265;
 wire clknet_1_0__leaf_net265;
 wire clknet_1_1__leaf_net265;
 wire clknet_0_net259;
 wire clknet_1_0__leaf_net259;
 wire clknet_1_1__leaf_net259;
 wire clknet_0_net691;
 wire clknet_1_0__leaf_net691;
 wire clknet_1_1__leaf_net691;
 wire clknet_0_net185;
 wire clknet_1_0__leaf_net185;
 wire clknet_1_1__leaf_net185;
 wire clknet_0_net868;
 wire clknet_1_0__leaf_net868;
 wire clknet_1_1__leaf_net868;
 wire clknet_0_net311;
 wire clknet_1_0__leaf_net311;
 wire clknet_1_1__leaf_net311;
 wire clknet_0_net287;
 wire clknet_1_0__leaf_net287;
 wire clknet_1_1__leaf_net287;
 wire clknet_0_net911;
 wire clknet_1_0__leaf_net911;
 wire clknet_1_1__leaf_net911;
 wire clknet_0_net306;
 wire clknet_1_0__leaf_net306;
 wire clknet_1_1__leaf_net306;
 wire clknet_0_net909;
 wire clknet_1_0__leaf_net909;
 wire clknet_1_1__leaf_net909;
 wire clknet_0_net307;
 wire clknet_1_0__leaf_net307;
 wire clknet_1_1__leaf_net307;
 wire clknet_0_net210;
 wire clknet_1_0__leaf_net210;
 wire clknet_1_1__leaf_net210;
 wire clknet_0_net187;
 wire clknet_1_0__leaf_net187;
 wire clknet_1_1__leaf_net187;
 wire clknet_0_net690;
 wire clknet_1_0__leaf_net690;
 wire clknet_1_1__leaf_net690;
 wire clknet_0_net880;
 wire clknet_1_0__leaf_net880;
 wire clknet_1_1__leaf_net880;
 wire clknet_0_net183;
 wire clknet_1_0__leaf_net183;
 wire clknet_1_1__leaf_net183;
 wire clknet_0_net689;
 wire clknet_1_0__leaf_net689;
 wire clknet_1_1__leaf_net689;
 wire clknet_0_net910;
 wire clknet_1_0__leaf_net910;
 wire clknet_1_1__leaf_net910;
 wire clknet_0_net673;
 wire clknet_1_0__leaf_net673;
 wire clknet_1_1__leaf_net673;
 wire clknet_0_net224;
 wire clknet_1_0__leaf_net224;
 wire clknet_1_1__leaf_net224;
 wire clknet_0_net649;
 wire clknet_1_0__leaf_net649;
 wire clknet_1_1__leaf_net649;
 wire clknet_0_net925;
 wire clknet_1_0__leaf_net925;
 wire clknet_1_1__leaf_net925;
 wire clknet_0_net304;
 wire clknet_1_0__leaf_net304;
 wire clknet_1_1__leaf_net304;
 wire clknet_0_net529;
 wire clknet_1_0__leaf_net529;
 wire clknet_1_1__leaf_net529;
 wire clknet_0_net202;
 wire clknet_1_0__leaf_net202;
 wire clknet_1_1__leaf_net202;
 wire clknet_0_net922;
 wire clknet_1_0__leaf_net922;
 wire clknet_1_1__leaf_net922;
 wire clknet_0_net100;
 wire clknet_1_0__leaf_net100;
 wire clknet_1_1__leaf_net100;
 wire clknet_0_net892;
 wire clknet_1_0__leaf_net892;
 wire clknet_1_1__leaf_net892;
 wire clknet_0_net672;
 wire clknet_1_0__leaf_net672;
 wire clknet_1_1__leaf_net672;
 wire clknet_0_net94;
 wire clknet_1_0__leaf_net94;
 wire clknet_1_1__leaf_net94;
 wire clknet_0_net325;
 wire clknet_1_0__leaf_net325;
 wire clknet_1_1__leaf_net325;
 wire clknet_0_net671;
 wire clknet_1_0__leaf_net671;
 wire clknet_1_1__leaf_net671;
 wire clknet_0_net88;
 wire clknet_1_0__leaf_net88;
 wire clknet_1_1__leaf_net88;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1068;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;

 sky130_fd_sc_hd__mux4_2 c100 (.A0(net855),
    .A1(net857),
    .A2(net852),
    .A3(net1032),
    .S0(net862),
    .S1(net833),
    .X(net0));
 sky130_fd_sc_hd__mux4_1 c101 (.A0(net849),
    .A1(net862),
    .A2(net857),
    .A3(net855),
    .S0(net856),
    .S1(net833),
    .X(net1));
 sky130_fd_sc_hd__mux4_2 c102 (.A0(net1028),
    .A1(net856),
    .A2(net857),
    .A3(net829),
    .S0(net847),
    .S1(net862),
    .X(net918));
 sky130_fd_sc_hd__mux4_2 c103 (.A0(net857),
    .A1(net849),
    .A2(net856),
    .A3(net862),
    .S0(net858),
    .S1(net815),
    .X(net938));
 sky130_fd_sc_hd__mux4_2 c104 (.A0(net1),
    .A1(net836),
    .A2(net852),
    .A3(net862),
    .S0(net848),
    .S1(net839),
    .X(net2));
 sky130_fd_sc_hd__mux4_2 c105 (.A0(net862),
    .A1(net857),
    .A2(net2),
    .A3(net856),
    .S0(net858),
    .S1(net1010),
    .X(net3));
 sky130_fd_sc_hd__mux4_1 c106 (.A0(net853),
    .A1(net858),
    .A2(net3),
    .A3(net836),
    .S0(net813),
    .S1(net1031),
    .X(net4));
 sky130_fd_sc_hd__mux4_2 c107 (.A0(net856),
    .A1(net4),
    .A2(net836),
    .A3(net855),
    .S0(net831),
    .S1(net862),
    .X(net905));
 sky130_fd_sc_hd__mux4_1 c108 (.A0(net2),
    .A1(net781),
    .A2(net863),
    .A3(net858),
    .S0(net835),
    .S1(net905),
    .X(net5));
 sky130_fd_sc_hd__mux4_2 c109 (.A0(net864),
    .A1(net836),
    .A2(net5),
    .A3(net3),
    .S0(net784),
    .S1(net905),
    .X(net920));
 sky130_fd_sc_hd__mux4_1 c110 (.A0(net1),
    .A1(net855),
    .A2(net818),
    .A3(net918),
    .S0(net815),
    .S1(net1017),
    .X(net6));
 sky130_fd_sc_hd__a41o_1 c111 (.A1(net790),
    .A2(net831),
    .A3(net819),
    .A4(net6),
    .B1(net1001),
    .X(net7));
 sky130_fd_sc_hd__a41o_1 c112 (.A1(net815),
    .A2(net842),
    .A3(net784),
    .A4(net1),
    .B1(net1017),
    .X(net8));
 sky130_fd_sc_hd__a41o_1 c113 (.A1(net853),
    .A2(net833),
    .A3(net847),
    .A4(net809),
    .B1(net819),
    .X(net916));
 sky130_fd_sc_hd__a41o_1 c114 (.A1(net8),
    .A2(net2),
    .A3(net809),
    .A4(net1001),
    .B1(net847),
    .X(net928));
 sky130_fd_sc_hd__mux4_1 c115 (.A0(net855),
    .A1(net831),
    .A2(net916),
    .A3(net858),
    .S0(net1017),
    .S1(net1001),
    .X(net937));
 sky130_fd_sc_hd__a41o_1 c116 (.A1(net784),
    .A2(net7),
    .A3(net938),
    .A4(net937),
    .B1(net787),
    .X(net927));
 sky130_fd_sc_hd__mux4_1 c117 (.A0(net844),
    .A1(net860),
    .A2(net8),
    .A3(net1004),
    .S0(net928),
    .S1(net818),
    .X(net9));
 sky130_fd_sc_hd__mux4_2 c118 (.A0(net833),
    .A1(net815),
    .A2(net937),
    .A3(net927),
    .S0(net1017),
    .S1(net8),
    .X(net10));
 sky130_fd_sc_hd__a41o_2 c119 (.A1(net1017),
    .A2(net10),
    .A3(net831),
    .A4(net1013),
    .B1(net818),
    .X(net11));
 sky130_fd_sc_hd__a41o_1 c120 (.A1(net784),
    .A2(net916),
    .A3(net1001),
    .A4(net818),
    .B1(net833),
    .X(net940));
 sky130_fd_sc_hd__a41o_1 c121 (.A1(net847),
    .A2(net11),
    .A3(net801),
    .A4(net844),
    .B1(net861),
    .X(net939));
 sky130_fd_sc_hd__a41o_1 c122 (.A1(net823),
    .A2(net812),
    .A3(net940),
    .A4(net809),
    .B1(net1017),
    .X(net930));
 sky130_fd_sc_hd__a41o_1 c123 (.A1(net6),
    .A2(net10),
    .A3(net930),
    .A4(net11),
    .B1(net940),
    .X(net941));
 sky130_fd_sc_hd__mux4_2 c124 (.A0(net1001),
    .A1(net784),
    .A2(net11),
    .A3(net818),
    .S0(net859),
    .S1(net1017),
    .X(net923));
 sky130_fd_sc_hd__mux4_2 c125 (.A0(net860),
    .A1(net862),
    .A2(net809),
    .A3(net842),
    .S0(net847),
    .S1(net784),
    .X(net914));
 sky130_fd_sc_hd__mux4_1 c126 (.A0(net9),
    .A1(net11),
    .A2(net817),
    .A3(net815),
    .S0(net839),
    .S1(net928),
    .X(net12));
 sky130_fd_sc_hd__mux4_1 c127 (.A0(net809),
    .A1(net930),
    .A2(net914),
    .A3(net847),
    .S0(net860),
    .S1(net941),
    .X(net886));
 sky130_fd_sc_hd__a41o_1 c128 (.A1(net12),
    .A2(net916),
    .A3(net930),
    .A4(net886),
    .B1(net853),
    .X(net942));
 sky130_fd_sc_hd__a41o_1 c129 (.A1(net842),
    .A2(net916),
    .A3(net914),
    .A4(net11),
    .B1(net819),
    .X(net13));
 sky130_fd_sc_hd__mux4_2 c130 (.A0(net13),
    .A1(net844),
    .A2(net942),
    .A3(net9),
    .S0(net10),
    .S1(net12),
    .X(net932));
 sky130_fd_sc_hd__mux4_1 c131 (.A0(net10),
    .A1(net914),
    .A2(net861),
    .A3(net905),
    .S0(net923),
    .S1(net932),
    .X(net14));
 sky130_fd_sc_hd__a41o_4 c132 (.A1(net1014),
    .A2(net1031),
    .A3(net1005),
    .A4(net1001),
    .B1(net1019),
    .X(net15));
 sky130_fd_sc_hd__a41o_4 c133 (.A1(net15),
    .A2(net999),
    .A3(net1030),
    .A4(net1000),
    .B1(net1028),
    .X(net16));
 sky130_fd_sc_hd__a31o_4 c134 (.A1(net999),
    .A2(net770),
    .A3(net1030),
    .B1(net1020),
    .X(net935));
 sky130_fd_sc_hd__a41o_4 c135 (.A1(net998),
    .A2(net1001),
    .A3(net770),
    .A4(net1031),
    .B1(net1004),
    .X(net17));
 sky130_fd_sc_hd__a41o_4 c136 (.A1(net17),
    .A2(net987),
    .A3(net1013),
    .A4(net1020),
    .B1(net1023),
    .X(net18));
 sky130_fd_sc_hd__a31o_4 c137 (.A1(net1006),
    .A2(net15),
    .A3(net1008),
    .B1(net1019),
    .X(net19));
 sky130_fd_sc_hd__a41o_4 c138 (.A1(net1000),
    .A2(net1030),
    .A3(net1010),
    .A4(net17),
    .B1(net987),
    .X(net865));
 sky130_fd_sc_hd__a41o_4 c139 (.A1(net987),
    .A2(net1001),
    .A3(net1012),
    .A4(net17),
    .B1(net986),
    .X(net20));
 sky130_fd_sc_hd__a41o_4 c140 (.A1(net1085),
    .A2(net1019),
    .A3(net1005),
    .A4(net982),
    .B1(net18),
    .X(net21));
 sky130_fd_sc_hd__a41o_4 c141 (.A1(net986),
    .A2(net1010),
    .A3(net1085),
    .A4(net1019),
    .B1(net978),
    .X(net22));
 sky130_fd_sc_hd__mux4_2 c142 (.A0(net22),
    .A1(net767),
    .A2(net1000),
    .A3(net982),
    .S0(net17),
    .S1(net1068),
    .X(net23));
 sky130_fd_sc_hd__a41o_4 c143 (.A1(net976),
    .A2(net767),
    .A3(net18),
    .A4(net982),
    .B1(net1068),
    .X(net24));
 sky130_fd_sc_hd__mux4_2 c144 (.A0(net976),
    .A1(net24),
    .A2(net1085),
    .A3(net982),
    .S0(net1019),
    .S1(net1068),
    .X(net25));
 sky130_fd_sc_hd__mux4_2 c145 (.A0(net982),
    .A1(net854),
    .A2(net25),
    .A3(net1085),
    .S0(net1033),
    .S1(net1030),
    .X(net26));
 sky130_fd_sc_hd__a41o_4 c146 (.A1(net26),
    .A2(net18),
    .A3(net1000),
    .A4(net978),
    .B1(net1049),
    .X(net27));
 sky130_fd_sc_hd__mux4_2 c147 (.A0(net17),
    .A1(net1030),
    .A2(net24),
    .A3(net987),
    .S0(net1019),
    .S1(net1068),
    .X(net28));
 sky130_fd_sc_hd__a41o_2 c148 (.A1(net975),
    .A2(net976),
    .A3(net25),
    .A4(net22),
    .B1(net1068),
    .X(net871));
 sky130_fd_sc_hd__a41o_4 c149 (.A1(net973),
    .A2(net22),
    .A3(net1068),
    .A4(net1085),
    .B1(net976),
    .X(net29));
 sky130_fd_sc_hd__mux4_2 c150 (.A0(net972),
    .A1(net767),
    .A2(net770),
    .A3(net987),
    .S0(net976),
    .S1(net973),
    .X(net30));
 sky130_fd_sc_hd__a41o_4 c151 (.A1(net1094),
    .A2(net975),
    .A3(net26),
    .A4(net971),
    .B1(net1068),
    .X(net881));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net1001),
    .A1(net969),
    .A2(net968),
    .A3(net1068),
    .S0(net1062),
    .S1(net971),
    .X(net31));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net964),
    .A1(net1038),
    .A2(net968),
    .A3(net22),
    .S0(net18),
    .S1(net975),
    .X(net32));
 sky130_fd_sc_hd__a41o_1 c154 (.A1(net792),
    .A2(net1023),
    .A3(net1024),
    .A4(net1004),
    .B1(net1020),
    .X(net33));
 sky130_fd_sc_hd__mux4_2 c155 (.A0(net1030),
    .A1(net33),
    .A2(net793),
    .A3(net1026),
    .S0(net1024),
    .S1(net792),
    .X(net34));
 sky130_fd_sc_hd__a41o_4 c156 (.A1(net18),
    .A2(net1002),
    .A3(net34),
    .A4(net973),
    .B1(net19),
    .X(net35));
 sky130_fd_sc_hd__mux4_2 c157 (.A0(net1062),
    .A1(net785),
    .A2(net786),
    .A3(net1026),
    .S0(net787),
    .S1(net1024),
    .X(net36));
 sky130_fd_sc_hd__a41o_1 c158 (.A1(net33),
    .A2(net22),
    .A3(net970),
    .A4(net973),
    .B1(net798),
    .X(net37));
 sky130_fd_sc_hd__a41o_2 c159 (.A1(net793),
    .A2(net999),
    .A3(net966),
    .A4(net1002),
    .B1(net36),
    .X(net38));
 sky130_fd_sc_hd__a41o_2 c160 (.A1(net1031),
    .A2(net1002),
    .A3(net36),
    .A4(net966),
    .B1(net970),
    .X(net913));
 sky130_fd_sc_hd__a41o_2 c161 (.A1(net963),
    .A2(net38),
    .A3(net33),
    .A4(net966),
    .B1(net970),
    .X(net39));
 sky130_fd_sc_hd__a41o_2 c162 (.A1(net1008),
    .A2(net793),
    .A3(net1006),
    .A4(net36),
    .B1(net33),
    .X(net924));
 sky130_fd_sc_hd__mux4_2 c163 (.A0(net770),
    .A1(net963),
    .A2(net1015),
    .A3(net786),
    .S0(net966),
    .S1(net970),
    .X(net40));
 sky130_fd_sc_hd__mux4_2 c164 (.A0(net959),
    .A1(net798),
    .A2(net1026),
    .A3(net971),
    .S0(net1028),
    .S1(net792),
    .X(net41));
 sky130_fd_sc_hd__mux4_2 c165 (.A0(net960),
    .A1(net924),
    .A2(net959),
    .A3(net767),
    .S0(net972),
    .S1(net1010),
    .X(net42));
 sky130_fd_sc_hd__a41o_2 c166 (.A1(net42),
    .A2(net770),
    .A3(net802),
    .A4(net999),
    .B1(net960),
    .X(net43));
 sky130_fd_sc_hd__a41o_1 c167 (.A1(net946),
    .A2(net785),
    .A3(net963),
    .A4(net966),
    .B1(net34),
    .X(net44));
 sky130_fd_sc_hd__mux4_2 c168 (.A0(net1006),
    .A1(net18),
    .A2(net959),
    .A3(net954),
    .S0(net924),
    .S1(net565),
    .X(net45));
 sky130_fd_sc_hd__mux4_1 c169 (.A0(net966),
    .A1(net45),
    .A2(net924),
    .A3(net33),
    .S0(net786),
    .S1(net1006),
    .X(net46));
 sky130_fd_sc_hd__mux4_2 c170 (.A0(net1031),
    .A1(net793),
    .A2(net780),
    .A3(net800),
    .S0(net785),
    .S1(net566),
    .X(net47));
 sky130_fd_sc_hd__mux4_2 c171 (.A0(net954),
    .A1(net794),
    .A2(net963),
    .A3(net47),
    .S0(net966),
    .S1(net959),
    .X(net48));
 sky130_fd_sc_hd__mux4_1 c172 (.A0(net38),
    .A1(net34),
    .A2(net960),
    .A3(net45),
    .S0(net47),
    .X(net49));
 sky130_fd_sc_hd__mux4_1 c173 (.A0(net786),
    .A1(net1013),
    .A2(net1100),
    .A3(net963),
    .S0(net48),
    .S1(net565),
    .X(net50));
 sky130_fd_sc_hd__a41o_1 c174 (.A1(net48),
    .A2(net38),
    .A3(net47),
    .A4(net1026),
    .B1(net566),
    .X(net51));
 sky130_fd_sc_hd__a41o_2 c175 (.A1(net47),
    .A2(net1031),
    .A3(net964),
    .A4(net566),
    .B1(net665),
    .X(net52));
 sky130_fd_sc_hd__mux4_2 c176 (.A0(net825),
    .A1(net820),
    .A2(net814),
    .A3(net18),
    .S0(net1005),
    .S1(net1028),
    .X(net53));
 sky130_fd_sc_hd__mux4_2 c177 (.A0(net18),
    .A1(net794),
    .A2(net924),
    .A3(net1024),
    .S0(net968),
    .S1(net664),
    .X(net54));
 sky130_fd_sc_hd__mux4_2 c178 (.A0(net816),
    .A1(net808),
    .A2(net1015),
    .A3(net805),
    .S0(net823),
    .S1(net817),
    .X(net55));
 sky130_fd_sc_hd__mux4_2 c179 (.A0(net1013),
    .A1(net814),
    .A2(net969),
    .A3(net822),
    .S0(net53),
    .S1(net1005),
    .X(net56));
 sky130_fd_sc_hd__a41o_1 c180 (.A1(net1026),
    .A2(net826),
    .A3(net804),
    .A4(net823),
    .B1(net1033),
    .X(net57));
 sky130_fd_sc_hd__a41o_4 c181 (.A1(net798),
    .A2(net57),
    .A3(net795),
    .A4(net54),
    .B1(net968),
    .X(net58));
 sky130_fd_sc_hd__a41o_2 c182 (.A1(net1023),
    .A2(net822),
    .A3(net827),
    .A4(net807),
    .B1(net1005),
    .X(net59));
 sky130_fd_sc_hd__mux4_2 c183 (.A0(net778),
    .A1(net825),
    .A2(net826),
    .A3(net814),
    .S0(net808),
    .S1(net816),
    .X(net884));
 sky130_fd_sc_hd__mux4_2 c184 (.A0(net785),
    .A1(net58),
    .A2(net963),
    .A3(net56),
    .S0(net57),
    .S1(net36),
    .X(net60));
 sky130_fd_sc_hd__a41o_2 c185 (.A1(net57),
    .A2(net55),
    .A3(net60),
    .A4(net54),
    .B1(net1015),
    .X(net61));
 sky130_fd_sc_hd__mux4_2 c186 (.A0(net807),
    .A1(net970),
    .A2(net56),
    .A3(net786),
    .S0(net53),
    .S1(net974),
    .X(net62));
 sky130_fd_sc_hd__mux4_2 c187 (.A0(net786),
    .A1(net56),
    .A2(net55),
    .A3(net812),
    .S0(net1032),
    .S1(net970),
    .X(net63));
 sky130_fd_sc_hd__mux4_2 c188 (.A0(net816),
    .A1(net1042),
    .A2(net56),
    .A3(net60),
    .S0(net798),
    .S1(net566),
    .X(net64));
 sky130_fd_sc_hd__mux4_1 c189 (.A0(net61),
    .A1(net806),
    .A2(net55),
    .A3(net60),
    .S0(net1005),
    .S1(net1043),
    .X(net65));
 sky130_fd_sc_hd__mux4_1 c190 (.A0(net59),
    .A1(net64),
    .A2(net55),
    .A3(net60),
    .S0(net1033),
    .S1(net579),
    .X(net66));
 sky130_fd_sc_hd__mux4_1 c191 (.A0(net884),
    .A1(net1016),
    .A2(net816),
    .A3(net946),
    .S0(net48),
    .X(net67));
 sky130_fd_sc_hd__mux4_1 c192 (.A0(net1042),
    .A1(net64),
    .A2(net978),
    .A3(net47),
    .S0(net816),
    .S1(net600),
    .X(net68));
 sky130_fd_sc_hd__mux4_1 c193 (.A0(net64),
    .A1(net823),
    .A2(net822),
    .A3(net827),
    .S0(net598),
    .S1(net600),
    .X(net69));
 sky130_fd_sc_hd__mux4_1 c194 (.A0(net807),
    .A1(net798),
    .A2(net45),
    .A3(net579),
    .S1(net667),
    .X(net70));
 sky130_fd_sc_hd__a41o_4 c195 (.A1(net978),
    .A2(net805),
    .A3(net59),
    .A4(net598),
    .B1(net666),
    .X(net71));
 sky130_fd_sc_hd__mux4_2 c196 (.A0(net60),
    .A1(net824),
    .A2(net54),
    .A3(net71),
    .S0(net598),
    .S1(net667),
    .X(net900));
 sky130_fd_sc_hd__mux4_1 c197 (.A0(net64),
    .A1(net794),
    .A2(net775),
    .S0(net598),
    .S1(net600),
    .X(net72));
 sky130_fd_sc_hd__mux4_1 c198 (.A0(net45),
    .A1(net830),
    .A2(net1016),
    .A3(net954),
    .S0(net61),
    .S1(net1018),
    .X(net73));
 sky130_fd_sc_hd__mux4_2 c199 (.A0(net1010),
    .A1(net831),
    .A2(net60),
    .A3(net959),
    .S0(net1051),
    .S1(net664),
    .X(net74));
 sky130_fd_sc_hd__mux4_1 c200 (.A0(net1050),
    .A1(net913),
    .A2(net54),
    .A3(net74),
    .S0(net850),
    .S1(net579),
    .X(net75));
 sky130_fd_sc_hd__mux4_1 c201 (.A0(net820),
    .A1(net833),
    .A2(net48),
    .A3(net1050),
    .S0(net877),
    .S1(net993),
    .X(net76));
 sky130_fd_sc_hd__mux4_1 c202 (.A0(net74),
    .A1(net813),
    .A2(net970),
    .A3(net820),
    .S0(net600),
    .S1(net993),
    .X(net77));
 sky130_fd_sc_hd__mux4_2 c203 (.A0(net1029),
    .A1(net59),
    .A2(net838),
    .A3(net1028),
    .S0(net1013),
    .S1(net995),
    .X(net78));
 sky130_fd_sc_hd__mux4_2 c204 (.A0(net840),
    .A1(net828),
    .A2(net781),
    .A3(net813),
    .S0(net993),
    .S1(net670),
    .X(net79));
 sky130_fd_sc_hd__mux4_2 c205 (.A0(net837),
    .A1(net78),
    .A2(net1015),
    .A3(net967),
    .S0(net664),
    .S1(net993),
    .X(net80));
 sky130_fd_sc_hd__mux4_2 c206 (.A0(net830),
    .A1(net78),
    .A2(net80),
    .A3(net1016),
    .S0(net840),
    .S1(net993),
    .X(net81));
 sky130_fd_sc_hd__mux4_2 c207 (.A0(net79),
    .A1(net78),
    .A2(net600),
    .A3(net994),
    .S0(net669),
    .S1(net670),
    .X(net82));
 sky130_fd_sc_hd__mux4_2 c208 (.A0(net785),
    .A1(net80),
    .A2(net82),
    .A3(net834),
    .S0(net1018),
    .S1(net993),
    .X(net83));
 sky130_fd_sc_hd__mux4_2 c209 (.A0(net81),
    .A1(net56),
    .A2(net82),
    .A3(net1033),
    .S0(net598),
    .S1(net993),
    .X(net84));
 sky130_fd_sc_hd__mux4_2 c210 (.A0(net835),
    .A1(net56),
    .A2(net81),
    .A3(net79),
    .S0(net578),
    .S1(net670),
    .X(net85));
 sky130_fd_sc_hd__mux4_1 c211 (.A0(net833),
    .A1(net1060),
    .A2(net61),
    .A3(net803),
    .S0(net598),
    .S1(net994),
    .X(net86));
 sky130_fd_sc_hd__mux4_2 c212 (.A0(net81),
    .A1(net953),
    .A2(net806),
    .A3(net851),
    .S0(net84),
    .S1(net1050),
    .X(net87));
 sky130_fd_sc_hd__mux4_1 c213 (.A0(net841),
    .A1(net34),
    .A2(net953),
    .A3(net812),
    .S0(net670),
    .S1(clknet_1_0__leaf_net671),
    .X(net88));
 sky130_fd_sc_hd__mux4_1 c214 (.A0(net824),
    .A1(net787),
    .A2(net80),
    .A3(net953),
    .S0(net898),
    .S1(net669),
    .X(net89));
 sky130_fd_sc_hd__mux4_1 c215 (.A0(net850),
    .A1(clknet_1_0__leaf_net88),
    .A2(net55),
    .A3(net953),
    .S0(net841),
    .S1(net578),
    .X(net90));
 sky130_fd_sc_hd__mux4_1 c216 (.A0(net827),
    .A1(net82),
    .A2(net89),
    .A3(net781),
    .S0(net578),
    .S1(net993),
    .X(net91));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(net83),
    .A1(net953),
    .A2(net1057),
    .A3(net781),
    .S0(clknet_1_0__leaf_net88),
    .X(net92));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(net55),
    .A1(net89),
    .A2(net82),
    .A3(net953),
    .S0(net592),
    .S1(net993),
    .X(net93));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net833),
    .A1(net15),
    .A2(net998),
    .A3(net592),
    .S0(net993),
    .S1(clknet_1_0__leaf_net672),
    .X(net94));
 sky130_fd_sc_hd__mux4_2 c220 (.A0(net1017),
    .A1(net84),
    .A2(net58),
    .A3(net839),
    .S0(net598),
    .S1(net994),
    .X(net929));
 sky130_fd_sc_hd__mux4_1 c221 (.A0(net48),
    .A1(net998),
    .A2(net3),
    .A3(net828),
    .S0(net1032),
    .S1(net665),
    .X(net95));
 sky130_fd_sc_hd__mux4_2 c222 (.A0(net829),
    .A1(net852),
    .A2(net998),
    .A3(net920),
    .S0(net857),
    .S1(net84),
    .X(net931));
 sky130_fd_sc_hd__mux4_2 c223 (.A0(net81),
    .A1(net0),
    .A2(net1008),
    .A3(net857),
    .S0(net1031),
    .S1(net972),
    .X(net96));
 sky130_fd_sc_hd__mux4_1 c224 (.A0(net961),
    .A1(net968),
    .A2(net831),
    .A3(net954),
    .S0(net87),
    .S1(net1031),
    .X(net97));
 sky130_fd_sc_hd__mux4_2 c225 (.A0(net781),
    .A1(net1028),
    .A2(net828),
    .A3(net938),
    .S0(net824),
    .S1(net675),
    .X(net98));
 sky130_fd_sc_hd__mux4_1 c226 (.A0(net62),
    .A1(net905),
    .A2(net45),
    .A3(net961),
    .S0(net790),
    .S1(net995),
    .X(net99));
 sky130_fd_sc_hd__mux4_1 c227 (.A0(net852),
    .A1(net1057),
    .A2(net963),
    .A3(net1013),
    .S0(net819),
    .S1(clknet_1_0__leaf_net673),
    .X(net100));
 sky130_fd_sc_hd__mux4_1 c228 (.A0(net848),
    .A1(net884),
    .A2(net1027),
    .A3(net920),
    .S0(net974),
    .S1(clknet_1_0__leaf_net673),
    .X(net922));
 sky130_fd_sc_hd__mux4_1 c229 (.A0(net87),
    .A1(clknet_1_1__leaf_net100),
    .A2(net1015),
    .A3(net848),
    .S0(net963),
    .S1(clknet_1_0__leaf_net673),
    .X(net101));
 sky130_fd_sc_hd__mux4_1 c230 (.A0(net87),
    .A1(net819),
    .A2(net963),
    .A3(clknet_1_0__leaf_net94),
    .S0(net62),
    .S1(clknet_1_0__leaf_net672),
    .X(net102));
 sky130_fd_sc_hd__mux4_1 c231 (.A0(net828),
    .A1(clknet_1_1__leaf_net100),
    .A2(net1028),
    .A3(net79),
    .S0(clknet_1_0__leaf_net672),
    .S1(net678),
    .X(net892));
 sky130_fd_sc_hd__mux4_1 c232 (.A0(net98),
    .A1(net58),
    .A2(net96),
    .A3(net53),
    .S0(net1017),
    .S1(net882),
    .X(net103));
 sky130_fd_sc_hd__mux4_2 c233 (.A0(net1031),
    .A1(net96),
    .A2(net938),
    .A3(net98),
    .S0(net882),
    .S1(net885),
    .X(net104));
 sky130_fd_sc_hd__mux4_1 c234 (.A0(clknet_1_0__leaf_net100),
    .A1(net104),
    .A2(net0),
    .A3(net839),
    .S0(net1017),
    .S1(net994),
    .X(net105));
 sky130_fd_sc_hd__mux4_1 c235 (.A0(net836),
    .A1(net104),
    .A2(net103),
    .A3(net87),
    .S0(net882),
    .S1(net678),
    .X(net106));
 sky130_fd_sc_hd__mux4_1 c236 (.A0(net98),
    .A1(net54),
    .A2(net835),
    .A3(net918),
    .S0(net901),
    .S1(net994),
    .X(net107));
 sky130_fd_sc_hd__mux4_1 c237 (.A0(net1042),
    .A1(net961),
    .A2(net1027),
    .A3(net592),
    .S0(net885),
    .S1(net679),
    .X(net108));
 sky130_fd_sc_hd__mux4_1 c238 (.A0(net84),
    .A1(net836),
    .A2(clknet_1_0__leaf_net892),
    .A3(net54),
    .S0(net104),
    .S1(net974),
    .X(net109));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net108),
    .A1(net79),
    .A2(net71),
    .A3(net864),
    .S0(net1031),
    .S1(net934),
    .X(net110));
 sky130_fd_sc_hd__mux4_1 c240 (.A0(net107),
    .A1(net108),
    .A2(net98),
    .A3(net839),
    .S0(net1024),
    .S1(net110),
    .X(net111));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(net5),
    .A1(net107),
    .A2(clknet_1_1__leaf_net922),
    .A3(net110),
    .S0(net882),
    .S1(net934),
    .X(net112));
 sky130_fd_sc_hd__mux4_1 c256 (.A0(net7),
    .A1(clknet_1_0__leaf_net100),
    .A2(net939),
    .A3(net1005),
    .S0(net920),
    .S1(net790),
    .X(net944));
 sky130_fd_sc_hd__mux4_2 c257 (.A0(net839),
    .A1(net11),
    .A2(net7),
    .A3(net916),
    .S0(net831),
    .S1(net934),
    .X(net113));
 sky130_fd_sc_hd__mux4_1 c258 (.A0(net113),
    .A1(net107),
    .A2(net920),
    .A3(net864),
    .S0(net932),
    .S1(net678),
    .X(net943));
 sky130_fd_sc_hd__mux4_1 c259 (.A0(net11),
    .A1(net931),
    .A2(net923),
    .A3(net113),
    .S0(net998),
    .S1(net934),
    .X(net114));
 sky130_fd_sc_hd__mux4_1 c260 (.A0(net110),
    .A1(net790),
    .A2(net839),
    .A3(net859),
    .S0(net938),
    .S1(net113),
    .X(net115));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(net823),
    .A1(net939),
    .A2(net113),
    .A3(net900),
    .S0(net933),
    .S1(net1080),
    .X(net116));
 sky130_fd_sc_hd__mux4_1 c262 (.A0(net53),
    .A1(net113),
    .A2(net858),
    .A3(net933),
    .S0(net915),
    .S1(net882),
    .X(net921));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net14),
    .A1(net864),
    .A2(net53),
    .A3(net800),
    .S0(net921),
    .S1(net915),
    .X(net945));
 sky130_fd_sc_hd__a41o_4 c264 (.A1(net1002),
    .A2(net24),
    .A3(net19),
    .A4(net1094),
    .B1(net1049),
    .X(net117));
 sky130_fd_sc_hd__a41o_4 c265 (.A1(net1012),
    .A2(net15),
    .A3(net998),
    .A4(net1018),
    .B1(net969),
    .X(net903));
 sky130_fd_sc_hd__a41o_1 c266 (.A1(net1023),
    .A2(net903),
    .A3(net1027),
    .A4(net23),
    .B1(net978),
    .X(net118));
 sky130_fd_sc_hd__a41o_2 c267 (.A1(net1014),
    .A2(net1034),
    .A3(net956),
    .A4(net778),
    .B1(net117),
    .X(net119));
 sky130_fd_sc_hd__a41o_4 c268 (.A1(net1000),
    .A2(net117),
    .A3(net1029),
    .A4(net956),
    .B1(net1103),
    .X(net120));
 sky130_fd_sc_hd__a41o_1 c269 (.A1(net117),
    .A2(net1040),
    .A3(net903),
    .A4(net955),
    .B1(net1000),
    .X(net121));
 sky130_fd_sc_hd__a41o_2 c270 (.A1(net120),
    .A2(net956),
    .A3(net1034),
    .A4(net117),
    .B1(net1006),
    .X(net122));
 sky130_fd_sc_hd__a41o_1 c271 (.A1(net1038),
    .A2(net117),
    .A3(net1062),
    .A4(net961),
    .B1(net955),
    .X(net123));
 sky130_fd_sc_hd__a41o_1 c272 (.A1(net1010),
    .A2(net121),
    .A3(net949),
    .A4(net22),
    .B1(net955),
    .X(net124));
 sky130_fd_sc_hd__a41o_1 c273 (.A1(net124),
    .A2(net119),
    .A3(net956),
    .A4(net950),
    .B1(net973),
    .X(net125));
 sky130_fd_sc_hd__mux4_1 c274 (.A0(net778),
    .A1(net122),
    .A2(net1068),
    .A3(net1027),
    .S0(net949),
    .S1(net955),
    .X(net126));
 sky130_fd_sc_hd__sdfbbn_2 c275 (.CLK_N(clknet_4_7_0_clk),
    .D(net770),
    .RESET_B(net949),
    .SCD(net122),
    .SCE(net955),
    .SET_B(net1071),
    .Q(net128),
    .Q_N(net127));
 sky130_fd_sc_hd__mux4_1 c276 (.A0(net1032),
    .A1(net124),
    .A2(net122),
    .A3(net1010),
    .S0(net949),
    .S1(net955),
    .X(net129));
 sky130_fd_sc_hd__a41o_1 c277 (.A1(net903),
    .A2(net121),
    .A3(net950),
    .A4(net955),
    .B1(net992),
    .X(net130));
 sky130_fd_sc_hd__a41o_2 c278 (.A1(net949),
    .A2(net1002),
    .A3(net955),
    .A4(net583),
    .B1(net590),
    .X(net131));
 sky130_fd_sc_hd__a41o_2 c279 (.A1(net1029),
    .A2(net128),
    .A3(net956),
    .A4(net1100),
    .B1(net949),
    .X(net132));
 sky130_fd_sc_hd__sdfbbn_2 c280 (.CLK_N(clknet_4_5_0_clk),
    .D(net767),
    .RESET_B(net949),
    .SCD(net122),
    .SCE(net955),
    .SET_B(net992),
    .Q(net134),
    .Q_N(net133));
 sky130_fd_sc_hd__mux4_1 c281 (.A0(net121),
    .A1(net130),
    .A2(net131),
    .A3(net949),
    .S0(net996),
    .S1(net1111),
    .X(net135));
 sky130_fd_sc_hd__mux4_2 c282 (.A0(net997),
    .A1(net1056),
    .A2(net950),
    .A3(net955),
    .S0(net583),
    .S1(net991),
    .X(net136));
 sky130_fd_sc_hd__mux4_1 c283 (.A0(net131),
    .A1(net121),
    .A2(net124),
    .A3(net996),
    .S0(net949),
    .S1(net991),
    .X(net137));
 sky130_fd_sc_hd__mux4_1 c284 (.A0(net122),
    .A1(net949),
    .A2(net997),
    .A3(net590),
    .S0(net992),
    .S1(net991),
    .X(net138));
 sky130_fd_sc_hd__mux4_1 c285 (.A0(net136),
    .A1(net997),
    .A2(net131),
    .A3(net767),
    .S0(net590),
    .S1(net990),
    .X(net139));
 sky130_fd_sc_hd__mux4_2 c286 (.A0(net768),
    .A1(net41),
    .A2(net1014),
    .A3(net959),
    .S0(net854),
    .S1(net565),
    .X(net140));
 sky130_fd_sc_hd__sdfbbp_1 c287 (.CLK(clknet_4_7_0_clk),
    .D(net803),
    .RESET_B(net997),
    .SCD(net132),
    .SCE(net41),
    .SET_B(net1077),
    .Q(net142),
    .Q_N(net141));
 sky130_fd_sc_hd__sdfbbn_2 c288 (.CLK_N(clknet_4_5_0_clk),
    .D(net33),
    .RESET_B(net951),
    .SCD(net27),
    .SCE(net946),
    .SET_B(net961),
    .Q(net144),
    .Q_N(net143));
 sky130_fd_sc_hd__a41o_1 c289 (.A1(net780),
    .A2(net144),
    .A3(net792),
    .A4(net664),
    .B1(net991),
    .X(net145));
 sky130_fd_sc_hd__mux4_2 c290 (.A0(net1015),
    .A1(net1030),
    .A2(net1111),
    .A3(net790),
    .S0(net780),
    .S1(net961),
    .X(net146));
 sky130_fd_sc_hd__sdfbbn_2 c291 (.CLK_N(clknet_4_4_0_clk),
    .D(net787),
    .RESET_B(net131),
    .SCD(net52),
    .SCE(net119),
    .SET_B(net1103),
    .Q(net148),
    .Q_N(net147));
 sky130_fd_sc_hd__mux4_2 c292 (.A0(net148),
    .A1(net801),
    .A2(net143),
    .A3(net1030),
    .S0(net117),
    .S1(net565),
    .X(net149));
 sky130_fd_sc_hd__a41o_1 c293 (.A1(net1056),
    .A2(net1030),
    .A3(net970),
    .A4(net1010),
    .B1(net1024),
    .X(net150));
 sky130_fd_sc_hd__mux4_1 c294 (.A0(net150),
    .A1(net146),
    .A2(net951),
    .A3(net946),
    .S0(net117),
    .S1(net991),
    .X(net151));
 sky130_fd_sc_hd__mux4_1 c295 (.A0(net130),
    .A1(net1015),
    .A2(net141),
    .A3(net147),
    .S0(net1068),
    .S1(net149),
    .X(net152));
 sky130_fd_sc_hd__a41o_4 c296 (.A1(net22),
    .A2(net966),
    .A3(net147),
    .A4(net780),
    .B1(net1067),
    .X(net153));
 sky130_fd_sc_hd__mux4_2 c297 (.A0(net971),
    .A1(net150),
    .A2(net36),
    .A3(net780),
    .S0(net924),
    .S1(net959),
    .X(net154));
 sky130_fd_sc_hd__mux4_2 c298 (.A0(net154),
    .A1(net52),
    .A2(net792),
    .A3(net145),
    .S0(net153),
    .S1(net978),
    .X(net155));
 sky130_fd_sc_hd__mux4_1 c299 (.A0(net132),
    .A1(net130),
    .A2(net154),
    .A3(net153),
    .S0(net155),
    .S1(net1081),
    .X(net156));
 sky130_fd_sc_hd__mux4_2 c300 (.A0(net145),
    .A1(net153),
    .A2(net154),
    .A3(net52),
    .S0(net1067),
    .S1(net685),
    .X(net157));
 sky130_fd_sc_hd__mux4_2 c301 (.A0(net34),
    .A1(net970),
    .A2(net153),
    .A3(net961),
    .S0(net974),
    .S1(net664),
    .X(net158));
 sky130_fd_sc_hd__mux4_1 c302 (.A0(net155),
    .A1(net145),
    .A2(net153),
    .A3(net770),
    .S0(net996),
    .S1(net1067),
    .X(net159));
 sky130_fd_sc_hd__sdfbbp_1 c303 (.CLK(clknet_4_5_0_clk),
    .D(net36),
    .RESET_B(net157),
    .SCD(net1035),
    .SCE(net153),
    .SET_B(net1073),
    .Q(net161),
    .Q_N(net160));
 sky130_fd_sc_hd__mux4_1 c304 (.A0(net161),
    .A1(net45),
    .A2(net913),
    .A3(net140),
    .S0(net877),
    .S1(net686),
    .X(net162));
 sky130_fd_sc_hd__mux4_2 c305 (.A0(net52),
    .A1(net153),
    .A2(net158),
    .A3(net778),
    .S0(net1081),
    .S1(net1084),
    .X(net163));
 sky130_fd_sc_hd__mux4_1 c306 (.A0(net163),
    .A1(net52),
    .A2(net140),
    .A3(net1072),
    .S0(net591),
    .S1(net992),
    .X(net164));
 sky130_fd_sc_hd__sdfbbn_1 c307 (.CLK_N(clknet_4_6_0_clk),
    .D(net121),
    .RESET_B(net153),
    .SCD(net132),
    .SCE(net158),
    .SET_B(net573),
    .Q(net166),
    .Q_N(net165));
 sky130_fd_sc_hd__mux4_2 c308 (.A0(net822),
    .A1(net42),
    .A2(net924),
    .A3(net1067),
    .S0(net991),
    .S1(net687),
    .X(net167));
 sky130_fd_sc_hd__mux4_2 c309 (.A0(net145),
    .A1(net999),
    .A2(net1016),
    .A3(net149),
    .S0(net120),
    .S1(net962),
    .X(net168));
 sky130_fd_sc_hd__a41o_2 c310 (.A1(net811),
    .A2(net161),
    .A3(net960),
    .A4(net999),
    .B1(net951),
    .X(net169));
 sky130_fd_sc_hd__a41o_1 c311 (.A1(net154),
    .A2(net822),
    .A3(net811),
    .A4(net167),
    .B1(net1083),
    .X(net170));
 sky130_fd_sc_hd__mux4_2 c312 (.A0(net150),
    .A1(net804),
    .A2(net768),
    .A3(net808),
    .S0(net959),
    .S1(net811),
    .X(net171));
 sky130_fd_sc_hd__mux4_1 c313 (.A0(net136),
    .A1(net171),
    .A2(net795),
    .A3(net42),
    .S0(net812),
    .S1(net1083),
    .X(net172));
 sky130_fd_sc_hd__mux4_1 c314 (.A0(net119),
    .A1(net813),
    .A2(net957),
    .A3(net884),
    .S0(net946),
    .S1(net167),
    .X(net173));
 sky130_fd_sc_hd__mux4_2 c315 (.A0(net986),
    .A1(net819),
    .A2(net171),
    .A3(net573),
    .S0(net877),
    .S1(net660),
    .X(net174));
 sky130_fd_sc_hd__mux4_1 c316 (.A0(net794),
    .A1(net169),
    .A2(net804),
    .A3(net167),
    .S0(net146),
    .S1(net42),
    .X(net175));
 sky130_fd_sc_hd__sdfbbn_2 c317 (.CLK_N(clknet_4_1_0_clk),
    .D(net167),
    .RESET_B(net168),
    .SCD(net960),
    .SCE(net1042),
    .SET_B(net899),
    .Q(net906),
    .Q_N(net176));
 sky130_fd_sc_hd__mux4_1 c318 (.A0(net64),
    .A1(net1028),
    .A2(net906),
    .A3(net168),
    .S0(net962),
    .S1(net171),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 c319 (.A0(net795),
    .A1(net174),
    .A2(net176),
    .A3(net962),
    .S0(net1045),
    .S1(net794),
    .X(net178));
 sky130_fd_sc_hd__mux4_1 c320 (.A0(net57),
    .A1(net906),
    .A2(net169),
    .A3(net122),
    .S0(net660),
    .S1(clknet_1_0__leaf_net689),
    .X(net179));
 sky130_fd_sc_hd__mux4_1 c321 (.A0(net174),
    .A1(net804),
    .A2(net171),
    .A3(net960),
    .S0(net659),
    .S1(clknet_1_0__leaf_net690),
    .X(net180));
 sky130_fd_sc_hd__mux4_1 c322 (.A0(net130),
    .A1(net167),
    .A2(net149),
    .A3(net822),
    .S0(clknet_1_0__leaf_net689),
    .S1(clknet_1_0__leaf_net691),
    .X(net181));
 sky130_fd_sc_hd__mux4_1 c323 (.A0(net787),
    .A1(net167),
    .A2(net168),
    .A3(net573),
    .S0(net594),
    .S1(clknet_1_0__leaf_net689),
    .X(net182));
 sky130_fd_sc_hd__mux4_1 c324 (.A0(net171),
    .A1(net954),
    .A2(clknet_1_0__leaf_net689),
    .A3(clknet_1_0__leaf_net690),
    .S0(net692),
    .S1(net694),
    .X(net183));
 sky130_fd_sc_hd__mux4_1 c325 (.A0(clknet_1_1__leaf_net183),
    .A1(net131),
    .A2(net169),
    .A3(net176),
    .S0(clknet_1_0__leaf_net689),
    .S1(clknet_1_0__leaf_net691),
    .X(net184));
 sky130_fd_sc_hd__mux4_1 c326 (.A0(net62),
    .A1(net903),
    .A2(net176),
    .A3(clknet_1_0__leaf_net691),
    .S0(net695),
    .S1(net893),
    .X(net185));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(net169),
    .A1(net130),
    .A2(clknet_1_0__leaf_net185),
    .A3(net1032),
    .S0(clknet_1_1__leaf_net183),
    .S1(net660),
    .X(net186));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(clknet_1_1__leaf_net185),
    .A1(net1013),
    .A2(net954),
    .A3(net659),
    .S0(clknet_1_0__leaf_net689),
    .S1(net696),
    .X(net187));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(clknet_1_0__leaf_net187),
    .A1(net146),
    .A2(clknet_1_0__leaf_net185),
    .A3(clknet_1_1__leaf_net183),
    .S0(net899),
    .S1(clknet_1_0__leaf_net689),
    .X(net188));
 sky130_fd_sc_hd__mux4_1 c330 (.A0(net89),
    .A1(net998),
    .A2(net813),
    .A3(net946),
    .S0(net1008),
    .S1(net787),
    .X(net189));
 sky130_fd_sc_hd__mux4_2 c331 (.A0(net838),
    .A1(net1100),
    .A2(net153),
    .A3(net974),
    .S0(net670),
    .S1(net694),
    .X(net190));
 sky130_fd_sc_hd__mux4_2 c332 (.A0(net153),
    .A1(net957),
    .A2(net1013),
    .A3(net790),
    .S0(net600),
    .S1(net695),
    .X(net191));
 sky130_fd_sc_hd__mux4_1 c333 (.A0(net60),
    .A1(net826),
    .A2(net919),
    .A3(net659),
    .S0(net899),
    .S1(net692),
    .X(net192));
 sky130_fd_sc_hd__mux4_1 c334 (.A0(net174),
    .A1(net85),
    .A2(net998),
    .A3(net143),
    .S0(net805),
    .S1(net919),
    .X(net193));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(net80),
    .A1(net1028),
    .A2(net163),
    .A3(net564),
    .S0(clknet_1_1__leaf_net911),
    .S1(net899),
    .X(net194));
 sky130_fd_sc_hd__mux4_1 c336 (.A0(net191),
    .A1(net954),
    .A2(net82),
    .A3(net995),
    .S0(clknet_1_0__leaf_net672),
    .S1(clknet_1_0__leaf_net689),
    .X(net910));
 sky130_fd_sc_hd__mux4_1 c337 (.A0(net192),
    .A1(net83),
    .A2(net845),
    .A3(net62),
    .S0(net578),
    .S1(clknet_1_0__leaf_net672),
    .X(net195));
 sky130_fd_sc_hd__mux4_2 c338 (.A0(net161),
    .A1(net935),
    .A2(net171),
    .A3(net696),
    .S0(net697),
    .S1(net698),
    .X(net196));
 sky130_fd_sc_hd__mux4_2 c339 (.A0(net834),
    .A1(net903),
    .A2(net817),
    .A3(net149),
    .S0(net697),
    .S1(net698),
    .X(net197));
 sky130_fd_sc_hd__mux4_1 c340 (.A0(net122),
    .A1(net191),
    .A2(net74),
    .A3(net1060),
    .S0(net197),
    .S1(net845),
    .X(net198));
 sky130_fd_sc_hd__mux4_2 c341 (.A0(net56),
    .A1(net42),
    .A2(net62),
    .A3(net1024),
    .S0(net626),
    .S1(net693),
    .X(net199));
 sky130_fd_sc_hd__mux4_2 c342 (.A0(net845),
    .A1(net835),
    .A2(net814),
    .A3(net953),
    .S0(net160),
    .S1(net191),
    .X(net888));
 sky130_fd_sc_hd__mux4_1 c343 (.A0(net163),
    .A1(net1012),
    .A2(net1045),
    .A3(net196),
    .S0(net659),
    .S1(net995),
    .X(net200));
 sky130_fd_sc_hd__mux4_1 c344 (.A0(net74),
    .A1(net196),
    .A2(net806),
    .A3(net967),
    .S0(net818),
    .S1(net698),
    .X(net201));
 sky130_fd_sc_hd__mux4_1 c345 (.A0(net149),
    .A1(net1001),
    .A2(net634),
    .A3(net902),
    .S0(clknet_1_1__leaf_net925),
    .S1(net919),
    .X(net202));
 sky130_fd_sc_hd__mux4_1 c346 (.A0(net971),
    .A1(clknet_1_0__leaf_net202),
    .A2(clknet_1_0__leaf_net185),
    .A3(net199),
    .S0(net963),
    .S1(net697),
    .X(net203));
 sky130_fd_sc_hd__mux4_1 c347 (.A0(clknet_1_0__leaf_net202),
    .A1(clknet_1_0__leaf_net183),
    .A2(net995),
    .A3(clknet_1_0__leaf_net689),
    .S0(net697),
    .S1(net904),
    .X(net204));
 sky130_fd_sc_hd__mux4_1 c348 (.A0(net851),
    .A1(clknet_1_1__leaf_net202),
    .A2(net171),
    .A3(net888),
    .S0(net662),
    .S1(net904),
    .X(net205));
 sky130_fd_sc_hd__mux4_1 c349 (.A0(clknet_1_1__leaf_net88),
    .A1(net199),
    .A2(net56),
    .A3(clknet_1_1__leaf_net911),
    .S0(net902),
    .S1(net697),
    .X(net206));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(clknet_1_1__leaf_net202),
    .A1(net199),
    .A2(net564),
    .A3(net626),
    .S0(net902),
    .S1(clknet_1_1__leaf_net925),
    .X(net207));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net192),
    .A1(net1082),
    .A2(net662),
    .A3(net995),
    .S0(net698),
    .S1(net1069),
    .X(net208));
 sky130_fd_sc_hd__mux4_1 c352 (.A0(net196),
    .A1(net859),
    .A2(net967),
    .A3(net1008),
    .S0(net803),
    .S1(net692),
    .X(net209));
 sky130_fd_sc_hd__mux4_1 c353 (.A0(net952),
    .A1(net148),
    .A2(net1042),
    .A3(net859),
    .S0(clknet_1_0__leaf_net911),
    .S1(clknet_1_1__leaf_net672),
    .X(net210));
 sky130_fd_sc_hd__mux4_1 c354 (.A0(clknet_1_0__leaf_net210),
    .A1(net972),
    .A2(net837),
    .A3(net888),
    .S0(net676),
    .S1(net695),
    .X(net211));
 sky130_fd_sc_hd__mux4_1 c355 (.A0(net813),
    .A1(net3),
    .A2(net98),
    .A3(net147),
    .S0(net837),
    .S1(net600),
    .X(net212));
 sky130_fd_sc_hd__mux4_1 c356 (.A0(net4),
    .A1(clknet_1_0__leaf_net210),
    .A2(net831),
    .A3(net212),
    .S0(net863),
    .S1(net882),
    .X(net213));
 sky130_fd_sc_hd__mux4_1 c357 (.A0(net0),
    .A1(net171),
    .A2(net826),
    .A3(net679),
    .S0(net899),
    .S1(net694),
    .X(net214));
 sky130_fd_sc_hd__mux4_1 c358 (.A0(net212),
    .A1(net931),
    .A2(net214),
    .A3(net1016),
    .S0(net835),
    .S1(net898),
    .X(net215));
 sky130_fd_sc_hd__mux4_1 c359 (.A0(net45),
    .A1(net920),
    .A2(net856),
    .A3(net635),
    .S0(net644),
    .S1(clknet_1_1__leaf_net672),
    .X(net216));
 sky130_fd_sc_hd__mux4_1 c360 (.A0(net214),
    .A1(net191),
    .A2(clknet_1_1__leaf_net910),
    .A3(net835),
    .S0(net3),
    .S1(net171),
    .X(net217));
 sky130_fd_sc_hd__mux4_1 c361 (.A0(net826),
    .A1(net801),
    .A2(net858),
    .A3(net831),
    .S0(net665),
    .S1(clknet_1_0__leaf_net671),
    .X(net917));
 sky130_fd_sc_hd__mux4_1 c362 (.A0(net863),
    .A1(net108),
    .A2(clknet_1_0__leaf_net892),
    .A3(net53),
    .S0(net859),
    .S1(net674),
    .X(net218));
 sky130_fd_sc_hd__mux4_1 c363 (.A0(net835),
    .A1(net214),
    .A2(clknet_1_0__leaf_net94),
    .A3(clknet_1_0__leaf_net925),
    .S0(net676),
    .S1(net904),
    .X(net219));
 sky130_fd_sc_hd__mux4_1 c364 (.A0(clknet_1_0__leaf_net910),
    .A1(net952),
    .A2(net627),
    .A3(clknet_1_1__leaf_net673),
    .S0(net684),
    .S1(net693),
    .X(net220));
 sky130_fd_sc_hd__mux4_1 c365 (.A0(net196),
    .A1(net929),
    .A2(net813),
    .A3(net1028),
    .S0(net644),
    .S1(clknet_1_0__leaf_net925),
    .X(net221));
 sky130_fd_sc_hd__mux4_1 c366 (.A0(net218),
    .A1(net171),
    .A2(net1032),
    .A3(net674),
    .S0(net697),
    .S1(net700),
    .X(net222));
 sky130_fd_sc_hd__mux4_1 c367 (.A0(net1042),
    .A1(net929),
    .A2(net199),
    .A3(net644),
    .S0(clknet_1_0__leaf_net671),
    .S1(net701),
    .X(net223));
 sky130_fd_sc_hd__mux4_1 c368 (.A0(net3),
    .A1(net191),
    .A2(net212),
    .A3(net906),
    .S0(net863),
    .S1(clknet_1_1__leaf_net673),
    .X(net224));
 sky130_fd_sc_hd__mux4_1 c369 (.A0(net824),
    .A1(clknet_1_0__leaf_net224),
    .A2(net635),
    .A3(net644),
    .S0(net675),
    .S1(net701),
    .X(net225));
 sky130_fd_sc_hd__mux4_1 c370 (.A0(net148),
    .A1(clknet_1_0__leaf_net224),
    .A2(net78),
    .A3(net627),
    .S0(net644),
    .S1(net701),
    .X(net226));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(clknet_1_0__leaf_net224),
    .A1(net600),
    .A2(net666),
    .A3(net670),
    .S0(clknet_1_1__leaf_net672),
    .S1(net701),
    .X(net227));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net58),
    .A1(clknet_1_1__leaf_net210),
    .A2(net1060),
    .A3(clknet_1_0__leaf_net224),
    .S0(clknet_1_0__leaf_net649),
    .S1(net697),
    .X(net228));
 sky130_fd_sc_hd__a41o_1 c373 (.A1(clknet_1_1__leaf_net224),
    .A2(net896),
    .A3(net644),
    .A4(clknet_1_0__leaf_net925),
    .B1(net662),
    .X(net229));
 sky130_fd_sc_hd__sdfbbp_1 c396 (.CLK(clknet_4_7_0_clk),
    .D(net124),
    .RESET_B(net1029),
    .SCD(net1061),
    .SCE(net973),
    .SET_B(net1000),
    .Q(net231),
    .Q_N(net230));
 sky130_fd_sc_hd__a41o_2 c397 (.A1(net969),
    .A2(net1010),
    .A3(net1014),
    .A4(net996),
    .B1(net979),
    .X(net232));
 sky130_fd_sc_hd__a41o_1 c398 (.A1(net231),
    .A2(net1051),
    .A3(net131),
    .A4(net1030),
    .B1(net590),
    .X(net233));
 sky130_fd_sc_hd__sdfbbn_2 c399 (.CLK_N(clknet_4_13_0_clk),
    .D(net1062),
    .RESET_B(net1051),
    .SCD(net1000),
    .SCE(net996),
    .SET_B(net136),
    .Q(net235),
    .Q_N(net234));
 sky130_fd_sc_hd__a41o_2 c400 (.A1(net231),
    .A2(net997),
    .A3(net1038),
    .A4(net776),
    .B1(net683),
    .X(net236));
 sky130_fd_sc_hd__a41o_2 c401 (.A1(net973),
    .A2(net24),
    .A3(net1012),
    .A4(net682),
    .B1(net683),
    .X(net237));
 sky130_fd_sc_hd__a41o_2 c402 (.A1(net237),
    .A2(net903),
    .A3(net1021),
    .A4(net964),
    .B1(net582),
    .X(net238));
 sky130_fd_sc_hd__mux4_2 c403 (.A0(net238),
    .A1(net767),
    .A2(net232),
    .A3(net582),
    .S0(net682),
    .S1(net683),
    .X(net239));
 sky130_fd_sc_hd__a41o_1 c404 (.A1(net235),
    .A2(net128),
    .A3(net1000),
    .A4(net119),
    .B1(net230),
    .X(net240));
 sky130_fd_sc_hd__a41o_2 c405 (.A1(net236),
    .A2(net1029),
    .A3(net232),
    .A4(net1012),
    .B1(net1000),
    .X(net241));
 sky130_fd_sc_hd__a41o_2 c406 (.A1(net237),
    .A2(net1034),
    .A3(net238),
    .A4(net935),
    .B1(net683),
    .X(net242));
 sky130_fd_sc_hd__sdfbbn_2 c407 (.CLK_N(clknet_4_7_0_clk),
    .D(net1056),
    .RESET_B(net241),
    .SCD(net240),
    .SCE(net236),
    .SET_B(net239),
    .Q(net244),
    .Q_N(net243));
 sky130_fd_sc_hd__a41o_4 c408 (.A1(net238),
    .A2(net239),
    .A3(net243),
    .A4(net996),
    .B1(net1021),
    .X(net245));
 sky130_fd_sc_hd__sdfbbp_1 c409 (.CLK(clknet_4_13_0_clk),
    .D(net240),
    .RESET_B(net241),
    .SCD(net973),
    .SCE(net230),
    .SET_B(net948),
    .Q(net247),
    .Q_N(net246));
 sky130_fd_sc_hd__mux4_1 c410 (.A0(net245),
    .A1(net768),
    .A2(net950),
    .A3(net956),
    .S0(net236),
    .S1(net582),
    .X(net248));
 sky130_fd_sc_hd__a41o_1 c411 (.A1(net244),
    .A2(net1062),
    .A3(net245),
    .A4(net238),
    .B1(net240),
    .X(net249));
 sky130_fd_sc_hd__mux4_2 c412 (.A0(net770),
    .A1(net237),
    .A2(net241),
    .A3(net997),
    .S0(net238),
    .S1(net703),
    .X(net250));
 sky130_fd_sc_hd__mux4_1 c413 (.A0(net124),
    .A1(net232),
    .A2(net243),
    .A3(net239),
    .S0(net854),
    .S1(net704),
    .X(net251));
 sky130_fd_sc_hd__mux4_1 c414 (.A0(net250),
    .A1(net16),
    .A2(net245),
    .A3(net582),
    .S0(net683),
    .S1(net703),
    .X(net252));
 sky130_fd_sc_hd__a41o_1 c415 (.A1(net241),
    .A2(net582),
    .A3(net703),
    .A4(net705),
    .B1(net706),
    .X(net253));
 sky130_fd_sc_hd__mux4_2 c416 (.A0(net1061),
    .A1(net948),
    .A2(net241),
    .A3(net246),
    .S0(net947),
    .S1(net706),
    .X(net254));
 sky130_fd_sc_hd__mux4_1 c417 (.A0(net254),
    .A1(net246),
    .A2(net230),
    .A3(net253),
    .S0(net704),
    .S1(net705),
    .X(net255));
 sky130_fd_sc_hd__mux4_2 c418 (.A0(net767),
    .A1(net165),
    .A2(net41),
    .A3(net34),
    .S0(net1032),
    .S1(net992),
    .X(net256));
 sky130_fd_sc_hd__mux4_2 c419 (.A0(net776),
    .A1(net146),
    .A2(net959),
    .A3(net34),
    .S0(net1111),
    .S1(net990),
    .X(net257));
 sky130_fd_sc_hd__mux4_1 c420 (.A0(net790),
    .A1(net237),
    .A2(net257),
    .A3(net254),
    .S0(net801),
    .S1(net992),
    .X(net258));
 sky130_fd_sc_hd__mux4_1 c421 (.A0(net146),
    .A1(net1056),
    .A2(net154),
    .A3(net1026),
    .S0(net582),
    .S1(clknet_1_1__leaf_net708),
    .X(net259));
 sky130_fd_sc_hd__sdfbbn_1 c422 (.CLK_N(clknet_4_6_0_clk),
    .D(net52),
    .RESET_B(net257),
    .SCD(net948),
    .SCE(net947),
    .SET_B(net801),
    .Q(net261),
    .Q_N(net260));
 sky130_fd_sc_hd__mux4_1 c423 (.A0(net1014),
    .A1(net997),
    .A2(net1073),
    .A3(net803),
    .S0(net800),
    .S1(clknet_1_1__leaf_net708),
    .X(net262));
 sky130_fd_sc_hd__sdfbbn_2 c424 (.CLK_N(clknet_4_7_0_clk),
    .D(net257),
    .RESET_B(clknet_1_0__leaf_net262),
    .SCD(net792),
    .SCE(net243),
    .SET_B(clknet_1_1__leaf_net708),
    .Q(net264),
    .Q_N(net263));
 sky130_fd_sc_hd__mux4_1 c425 (.A0(net117),
    .A1(net166),
    .A2(net263),
    .A3(net999),
    .S0(clknet_1_0__leaf_net262),
    .S1(net800),
    .X(net265));
 sky130_fd_sc_hd__mux4_1 c426 (.A0(net254),
    .A1(net261),
    .A2(net237),
    .A3(net52),
    .S0(net257),
    .S1(net801),
    .X(net266));
 sky130_fd_sc_hd__sdfbbp_1 c427 (.CLK(clknet_4_7_0_clk),
    .D(clknet_1_1__leaf_net262),
    .RESET_B(net256),
    .SCD(net165),
    .SCE(net1061),
    .SET_B(net854),
    .Q(net268),
    .Q_N(net267));
 sky130_fd_sc_hd__sdfbbn_1 c428 (.CLK_N(clknet_4_12_0_clk),
    .D(net1016),
    .RESET_B(net16),
    .SCD(net257),
    .SCE(net267),
    .SET_B(net1036),
    .Q(net270),
    .Q_N(net269));
 sky130_fd_sc_hd__mux4_2 c429 (.A0(net795),
    .A1(net38),
    .A2(net260),
    .A3(net234),
    .S0(net573),
    .S1(net580),
    .X(net271));
 sky130_fd_sc_hd__a41o_2 c430 (.A1(net1085),
    .A2(net263),
    .A3(net271),
    .A4(net1024),
    .B1(net582),
    .X(net272));
 sky130_fd_sc_hd__mux4_1 c431 (.A0(clknet_1_1__leaf_net259),
    .A1(net35),
    .A2(net256),
    .A3(net264),
    .S0(net272),
    .S1(clknet_1_1__leaf_net708),
    .X(net273));
 sky130_fd_sc_hd__mux4_1 c432 (.A0(clknet_1_0__leaf_net265),
    .A1(net35),
    .A2(clknet_1_1__leaf_net259),
    .A3(net232),
    .S0(net269),
    .S1(net705),
    .X(net274));
 sky130_fd_sc_hd__mux4_1 c433 (.A0(net272),
    .A1(net267),
    .A2(net966),
    .A3(net1021),
    .S0(net580),
    .S1(clknet_1_0__leaf_net709),
    .X(net275));
 sky130_fd_sc_hd__mux4_1 c434 (.A0(net999),
    .A1(clknet_1_0__leaf_net275),
    .A2(net271),
    .A3(clknet_1_1__leaf_net265),
    .S0(clknet_1_1__leaf_net259),
    .S1(net36),
    .X(net276));
 sky130_fd_sc_hd__a41o_1 c435 (.A1(net957),
    .A2(net272),
    .A3(net947),
    .A4(net573),
    .B1(clknet_1_1__leaf_net875),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net270),
    .A1(clknet_1_1__leaf_net265),
    .A2(net263),
    .A3(net580),
    .S0(net594),
    .S1(clknet_1_1__leaf_net875),
    .X(net278));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(clknet_1_1__leaf_net277),
    .A1(clknet_1_0__leaf_net265),
    .A2(clknet_1_0__leaf_net278),
    .A3(net1033),
    .S0(net960),
    .S1(clknet_1_1__leaf_net875),
    .X(net279));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(clknet_1_1__leaf_net259),
    .A1(net272),
    .A2(clknet_1_1__leaf_net277),
    .A3(net263),
    .S0(clknet_1_0__leaf_net709),
    .S1(clknet_1_1__leaf_net875),
    .X(net280));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net261),
    .A1(clknet_1_1__leaf_net277),
    .A2(net166),
    .A3(clknet_1_0__leaf_net278),
    .S1(net619),
    .X(net281));
 sky130_fd_sc_hd__mux4_1 c440 (.A0(net1016),
    .A1(net168),
    .A2(net58),
    .A3(clknet_1_1__leaf_net277),
    .S0(net1029),
    .S1(net157),
    .X(net282));
 sky130_fd_sc_hd__mux4_1 c441 (.A0(net131),
    .A1(net900),
    .A2(net1060),
    .A3(net154),
    .S0(clknet_1_1__leaf_net875),
    .S1(net710),
    .X(net283));
 sky130_fd_sc_hd__mux4_1 c442 (.A0(net169),
    .A1(net803),
    .A2(net974),
    .A3(net999),
    .S0(net591),
    .S1(net683),
    .X(net284));
 sky130_fd_sc_hd__mux4_1 c443 (.A0(clknet_1_1__leaf_net187),
    .A1(net247),
    .A2(clknet_1_0__leaf_net277),
    .A3(net245),
    .S0(clknet_1_1__leaf_net689),
    .S1(net712),
    .X(net285));
 sky130_fd_sc_hd__mux4_2 c444 (.A0(net1012),
    .A1(net808),
    .A2(net975),
    .A3(net710),
    .S0(net712),
    .S1(net714),
    .X(net286));
 sky130_fd_sc_hd__mux4_1 c445 (.A0(net804),
    .A1(net812),
    .A2(net824),
    .A3(clknet_1_0__leaf_net185),
    .S0(net286),
    .S1(net959),
    .X(net287));
 sky130_fd_sc_hd__mux4_1 c446 (.A0(net158),
    .A1(net1006),
    .A2(net286),
    .A3(net27),
    .S0(net615),
    .S1(net714),
    .X(net288));
 sky130_fd_sc_hd__mux4_1 c447 (.A0(net168),
    .A1(net802),
    .A2(clknet_1_0__leaf_net259),
    .A3(net286),
    .S0(net619),
    .S1(net711),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 c448 (.A0(net168),
    .A1(net260),
    .A2(net47),
    .A3(net615),
    .S0(clknet_1_1__leaf_net690),
    .S1(clknet_1_0__leaf_net709),
    .X(net290));
 sky130_fd_sc_hd__mux4_1 c449 (.A0(net999),
    .A1(net957),
    .A2(net806),
    .A3(net992),
    .S0(net688),
    .S1(net908),
    .X(net291));
 sky130_fd_sc_hd__mux4_1 c450 (.A0(net62),
    .A1(net975),
    .A2(net237),
    .A3(net291),
    .S0(net1015),
    .S1(net688),
    .X(net292));
 sky130_fd_sc_hd__mux4_2 c451 (.A0(net997),
    .A1(net800),
    .A2(clknet_1_0__leaf_net278),
    .A3(net1050),
    .S0(net713),
    .S1(net716),
    .X(net293));
 sky130_fd_sc_hd__mux4_1 c452 (.A0(clknet_1_0__leaf_net287),
    .A1(net47),
    .A2(net58),
    .A3(net978),
    .S0(net168),
    .S1(net715),
    .X(net294));
 sky130_fd_sc_hd__mux4_1 c453 (.A0(net292),
    .A1(clknet_1_0__leaf_net277),
    .A2(net256),
    .A3(net991),
    .S0(clknet_1_0__leaf_net690),
    .S1(net717),
    .X(net295));
 sky130_fd_sc_hd__mux4_1 c454 (.A0(net142),
    .A1(net40),
    .A2(clknet_1_0__leaf_net293),
    .A3(net948),
    .S0(net615),
    .S1(net717),
    .X(net912));
 sky130_fd_sc_hd__mux4_2 c455 (.A0(net247),
    .A1(net618),
    .A2(net647),
    .A3(net660),
    .S0(net908),
    .S1(net717),
    .X(net296));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(net291),
    .A1(net292),
    .A2(clknet_1_0__leaf_net293),
    .A3(clknet_1_1__leaf_net912),
    .S0(net647),
    .S1(net713),
    .X(net297));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(net288),
    .A1(clknet_1_1__leaf_net912),
    .A2(clknet_1_0__leaf_net275),
    .A3(net615),
    .S0(net647),
    .S1(net718),
    .X(net298));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(net806),
    .A1(net795),
    .A2(net966),
    .A3(net36),
    .S0(net710),
    .S1(net718),
    .X(net299));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net947),
    .A1(clknet_1_0__leaf_net278),
    .A2(net615),
    .A3(net618),
    .S0(net666),
    .S1(net715),
    .X(net300));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net299),
    .A1(net174),
    .A2(net296),
    .A3(net168),
    .S0(net269),
    .S1(net990),
    .X(net301));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net299),
    .A1(net168),
    .A2(clknet_1_0__leaf_net278),
    .A3(net618),
    .S0(clknet_1_1__leaf_net689),
    .S1(net988),
    .X(net302));
 sky130_fd_sc_hd__mux4_1 c462 (.A0(net806),
    .A1(net244),
    .A2(clknet_1_0__leaf_net293),
    .A3(net42),
    .S0(net967),
    .S1(net662),
    .X(net303));
 sky130_fd_sc_hd__mux4_2 c463 (.A0(net837),
    .A1(net244),
    .A2(net964),
    .A3(clknet_1_1__leaf_net925),
    .S0(net698),
    .S1(net908),
    .X(net304));
 sky130_fd_sc_hd__mux4_1 c464 (.A0(net82),
    .A1(clknet_1_1__leaf_net910),
    .A2(clknet_1_0__leaf_net303),
    .A3(net190),
    .S0(net584),
    .S1(net908),
    .X(net305));
 sky130_fd_sc_hd__mux4_1 c465 (.A0(net971),
    .A1(net1003),
    .A2(clknet_1_1__leaf_net911),
    .A3(net648),
    .S0(net698),
    .S1(net716),
    .X(net306));
 sky130_fd_sc_hd__mux4_1 c466 (.A0(net947),
    .A1(clknet_1_0__leaf_net306),
    .A2(net1057),
    .A3(net669),
    .S0(net688),
    .S1(net716),
    .X(net307));
 sky130_fd_sc_hd__mux4_1 c467 (.A0(clknet_1_1__leaf_net303),
    .A1(net1008),
    .A2(net947),
    .A3(net174),
    .S0(net600),
    .S1(clknet_1_1__leaf_net672),
    .X(net308));
 sky130_fd_sc_hd__mux4_1 c468 (.A0(net174),
    .A1(clknet_1_0__leaf_net307),
    .A2(net947),
    .A3(net264),
    .S0(net1013),
    .S1(net635),
    .X(net309));
 sky130_fd_sc_hd__mux4_1 c469 (.A0(net237),
    .A1(clknet_1_1__leaf_net307),
    .A2(net806),
    .A3(clknet_1_1__leaf_net911),
    .S0(net688),
    .S1(net720),
    .X(net310));
 sky130_fd_sc_hd__mux4_1 c470 (.A0(clknet_1_1__leaf_net185),
    .A1(net1005),
    .A2(net574),
    .A3(net622),
    .S0(net904),
    .S1(net721),
    .X(net311));
 sky130_fd_sc_hd__mux4_1 c471 (.A0(clknet_1_1__leaf_net307),
    .A1(net158),
    .A2(net838),
    .A3(net1027),
    .S0(net71),
    .S1(net1082),
    .X(net312));
 sky130_fd_sc_hd__mux4_2 c472 (.A0(net15),
    .A1(net837),
    .A2(net954),
    .A3(net234),
    .S0(net564),
    .S1(net995),
    .X(net872));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(clknet_1_1__leaf_net185),
    .A1(net231),
    .A2(net1008),
    .A3(net574),
    .S0(net621),
    .S1(net988),
    .X(net868));
 sky130_fd_sc_hd__mux4_1 c474 (.A0(clknet_1_0__leaf_net307),
    .A1(net806),
    .A2(net54),
    .A3(net626),
    .S0(clknet_1_0__leaf_net708),
    .S1(net721),
    .X(net313));
 sky130_fd_sc_hd__mux4_2 c475 (.A0(clknet_1_0__leaf_net304),
    .A1(clknet_1_0__leaf_net293),
    .A2(net53),
    .A3(net817),
    .S0(net574),
    .S1(net662),
    .X(net314));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(net1050),
    .A1(clknet_1_0__leaf_net307),
    .A2(net837),
    .A3(net584),
    .S0(net634),
    .S1(clknet_1_1__leaf_net925),
    .X(net315));
 sky130_fd_sc_hd__mux4_2 c477 (.A0(net59),
    .A1(clknet_1_0__leaf_net304),
    .A2(net296),
    .A3(clknet_1_1__leaf_net314),
    .S0(net622),
    .S1(net883),
    .X(net316));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(net888),
    .A1(net1087),
    .A2(clknet_1_0__leaf_net311),
    .A3(clknet_1_0__leaf_net316),
    .S0(net574),
    .S1(clknet_1_0__leaf_net911),
    .X(net317));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(clknet_1_1__leaf_net311),
    .A1(clknet_1_0__leaf_net868),
    .A2(net83),
    .A3(net897),
    .S0(net669),
    .S1(clknet_1_0__leaf_net671),
    .X(net318));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(clknet_1_0__leaf_net304),
    .A1(net144),
    .A2(clknet_1_0__leaf_net306),
    .A3(net646),
    .S0(net656),
    .S1(net716),
    .X(net909));
 sky130_fd_sc_hd__mux4_2 c481 (.A0(net1094),
    .A1(net120),
    .A2(net35),
    .A3(net646),
    .S0(net656),
    .S1(net723),
    .X(net319));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(net231),
    .A1(net319),
    .A2(net656),
    .A3(net720),
    .S0(net722),
    .S1(net723),
    .X(net320));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(clknet_1_0__leaf_net314),
    .A1(net1087),
    .A2(net319),
    .A3(clknet_1_0__leaf_net311),
    .S0(net1008),
    .S1(net655),
    .X(net321));
 sky130_fd_sc_hd__mux4_1 c484 (.A0(net103),
    .A1(clknet_1_0__leaf_net183),
    .A2(net1018),
    .A3(net78),
    .S0(net859),
    .S1(net905),
    .X(net322));
 sky130_fd_sc_hd__mux4_1 c485 (.A0(net856),
    .A1(clknet_1_1__leaf_net94),
    .A2(clknet_1_1__leaf_net224),
    .A3(net837),
    .S0(net675),
    .S1(clknet_1_0__leaf_net708),
    .X(net323));
 sky130_fd_sc_hd__mux4_1 c486 (.A0(net96),
    .A1(net98),
    .A2(net199),
    .A3(net1013),
    .S0(net915),
    .S1(net662),
    .X(net324));
 sky130_fd_sc_hd__mux4_1 c487 (.A0(clknet_1_1__leaf_net94),
    .A1(net801),
    .A2(net817),
    .A3(net1003),
    .S0(net670),
    .S1(net702),
    .X(net325));
 sky130_fd_sc_hd__mux4_1 c488 (.A0(net104),
    .A1(clknet_1_0__leaf_net912),
    .A2(net96),
    .A3(clknet_1_0__leaf_net894),
    .S0(net628),
    .S1(net702),
    .X(net326));
 sky130_fd_sc_hd__mux4_1 c489 (.A0(net1014),
    .A1(net655),
    .A2(net662),
    .A3(net670),
    .S0(net678),
    .S1(net679),
    .X(net327));
 sky130_fd_sc_hd__mux4_2 c490 (.A0(net98),
    .A1(net1008),
    .A2(net972),
    .A3(net902),
    .S0(net685),
    .S1(net693),
    .X(net328));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(net261),
    .A1(net319),
    .A2(net327),
    .A3(net628),
    .S0(net655),
    .S1(net684),
    .X(net329));
 sky130_fd_sc_hd__mux4_1 c492 (.A0(net857),
    .A1(net952),
    .A2(net948),
    .A3(net328),
    .S0(clknet_1_1__leaf_net894),
    .S1(net679),
    .X(net330));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(net268),
    .A1(clknet_1_1__leaf_net224),
    .A2(net797),
    .A3(net594),
    .S0(net677),
    .S1(net685),
    .X(net331));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(net96),
    .A1(net328),
    .A2(net158),
    .A3(net594),
    .S0(net626),
    .S1(clknet_1_1__leaf_net672),
    .X(net895));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(net961),
    .A1(net856),
    .A2(net896),
    .A3(net625),
    .S0(net679),
    .S1(net717),
    .X(net332));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(net158),
    .A1(net257),
    .A2(net332),
    .A3(net901),
    .S0(net902),
    .S1(net701),
    .X(net333));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net327),
    .A1(clknet_1_0__leaf_net293),
    .A2(net594),
    .A3(net598),
    .S0(clknet_1_1__leaf_net672),
    .S1(net702),
    .X(net334));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(net846),
    .A1(net625),
    .A2(net700),
    .A3(clknet_1_0__leaf_net708),
    .S0(net883),
    .S1(net723),
    .X(net335));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(clknet_1_0__leaf_net335),
    .A1(net918),
    .A2(net946),
    .A3(net819),
    .S0(net877),
    .S1(clknet_1_1__leaf_net894),
    .X(net336));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(net334),
    .A1(net142),
    .A2(net837),
    .A3(clknet_1_1__leaf_net224),
    .S0(clknet_1_1__leaf_net335),
    .S1(net1085),
    .X(net337));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(net837),
    .A1(clknet_1_0__leaf_net335),
    .A2(net856),
    .A3(net901),
    .S0(net995),
    .S1(net686),
    .X(net907));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(net78),
    .A1(net833),
    .A2(clknet_1_0__leaf_net907),
    .A3(net1007),
    .S0(net1027),
    .S1(net677),
    .X(net338));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(net1060),
    .A1(net332),
    .A2(clknet_1_1__leaf_net907),
    .A3(clknet_1_1__leaf_net892),
    .S0(net857),
    .S1(net988),
    .X(net339));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net199),
    .A1(net244),
    .A2(net120),
    .A3(net332),
    .S0(clknet_1_1__leaf_net907),
    .S1(net662),
    .X(net340));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(clknet_1_0__leaf_net330),
    .A1(net53),
    .A2(net268),
    .A3(clknet_1_0__leaf_net338),
    .S0(clknet_1_1__leaf_net907),
    .S1(net1080),
    .X(net341));
 sky130_fd_sc_hd__a41o_4 c528 (.A1(net250),
    .A2(net1045),
    .A3(net239),
    .A4(net971),
    .B1(net1021),
    .X(net342));
 sky130_fd_sc_hd__a41o_1 c529 (.A1(net232),
    .A2(net968),
    .A3(net981),
    .A4(net958),
    .B1(net584),
    .X(net343));
 sky130_fd_sc_hd__a41o_1 c530 (.A1(net132),
    .A2(net958),
    .A3(net1006),
    .A4(net236),
    .B1(net1076),
    .X(net344));
 sky130_fd_sc_hd__mux4_1 c531 (.A0(net240),
    .A1(net247),
    .A2(net1003),
    .A3(net948),
    .S0(net1021),
    .S1(net705),
    .X(net345));
 sky130_fd_sc_hd__a41o_2 c532 (.A1(net119),
    .A2(net1038),
    .A3(net962),
    .A4(net236),
    .B1(net1105),
    .X(net346));
 sky130_fd_sc_hd__a41o_2 c533 (.A1(net1033),
    .A2(net343),
    .A3(net1051),
    .A4(net996),
    .B1(net1061),
    .X(net889));
 sky130_fd_sc_hd__sdfbbn_1 c534 (.CLK_N(clknet_4_13_0_clk),
    .D(net973),
    .RESET_B(net343),
    .SCD(net346),
    .SCE(net238),
    .SET_B(net704),
    .Q(net348),
    .Q_N(net347));
 sky130_fd_sc_hd__a41o_4 c535 (.A1(net241),
    .A2(net250),
    .A3(net1010),
    .A4(net1021),
    .B1(net724),
    .X(net349));
 sky130_fd_sc_hd__mux4_1 c536 (.A0(net889),
    .A1(net349),
    .A2(net346),
    .A3(net1054),
    .S0(net1021),
    .S1(net582),
    .X(net350));
 sky130_fd_sc_hd__mux4_1 c537 (.A0(net773),
    .A1(net349),
    .A2(net1054),
    .A3(net1021),
    .S0(net568),
    .S1(net705),
    .X(net351));
 sky130_fd_sc_hd__sdfbbp_1 c538 (.CLK(clknet_4_15_0_clk),
    .D(net343),
    .RESET_B(net349),
    .SCD(net1006),
    .SCE(net342),
    .SET_B(net1070),
    .Q(net353),
    .Q_N(net352));
 sky130_fd_sc_hd__sdfbbn_1 c539 (.CLK_N(clknet_4_15_0_clk),
    .D(net349),
    .RESET_B(net958),
    .SCD(net971),
    .SCE(net1014),
    .SET_B(net352),
    .Q(net355),
    .Q_N(net354));
 sky130_fd_sc_hd__mux4_1 c540 (.A0(net342),
    .A1(net346),
    .A2(net1011),
    .A3(net1012),
    .S0(net250),
    .S1(net1061),
    .X(net356));
 sky130_fd_sc_hd__mux4_2 c541 (.A0(net25),
    .A1(net1029),
    .A2(net347),
    .A3(net583),
    .S0(net707),
    .S1(net725),
    .X(net357));
 sky130_fd_sc_hd__sdfbbn_1 c542 (.CLK_N(clknet_4_13_0_clk),
    .D(net1027),
    .RESET_B(net881),
    .SCD(net240),
    .SCE(net706),
    .SET_B(clknet_1_1__leaf_net726),
    .Q(net359),
    .Q_N(net358));
 sky130_fd_sc_hd__mux4_1 c543 (.A0(net353),
    .A1(net342),
    .A2(net1048),
    .A3(net1057),
    .S0(net358),
    .S1(net250),
    .X(net360));
 sky130_fd_sc_hd__a41o_1 c544 (.A1(net348),
    .A2(net354),
    .A3(net584),
    .A4(clknet_1_1__leaf_net726),
    .B1(clknet_1_1__leaf_net727),
    .X(net361));
 sky130_fd_sc_hd__mux4_1 c545 (.A0(net236),
    .A1(net1006),
    .A2(net346),
    .A3(net240),
    .S0(clknet_1_1__leaf_net361),
    .S1(clknet_1_1__leaf_net727),
    .X(net362));
 sky130_fd_sc_hd__a41o_1 c546 (.A1(net128),
    .A2(net359),
    .A3(clknet_1_0__leaf_net361),
    .A4(net357),
    .B1(clknet_1_1__leaf_net727),
    .X(net363));
 sky130_fd_sc_hd__a41o_1 c547 (.A1(net979),
    .A2(net1033),
    .A3(net354),
    .A4(clknet_1_0__leaf_net363),
    .B1(clknet_1_1__leaf_net727),
    .X(net364));
 sky130_fd_sc_hd__mux4_1 c548 (.A0(net238),
    .A1(clknet_1_0__leaf_net363),
    .A2(net355),
    .A3(net1023),
    .S0(clknet_1_1__leaf_net727),
    .S1(clknet_1_1__leaf_net728),
    .X(net365));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(net239),
    .A1(clknet_1_1__leaf_net361),
    .A2(clknet_1_1__leaf_net363),
    .A3(net346),
    .S0(net951),
    .S1(net568),
    .X(net366));
 sky130_fd_sc_hd__mux4_1 c550 (.A0(net166),
    .A1(net348),
    .A2(net1027),
    .A3(net246),
    .S0(net263),
    .S1(net1026),
    .X(net869));
 sky130_fd_sc_hd__mux4_1 c551 (.A0(net140),
    .A1(net984),
    .A2(net232),
    .A3(net263),
    .S0(net683),
    .S1(clknet_1_1__leaf_net727),
    .X(net367));
 sky130_fd_sc_hd__mux4_1 c552 (.A0(net142),
    .A1(net165),
    .A2(net986),
    .A3(net234),
    .S0(net962),
    .S1(clknet_1_1__leaf_net727),
    .X(net368));
 sky130_fd_sc_hd__mux4_1 c553 (.A0(clknet_1_0__leaf_net368),
    .A1(net1037),
    .A2(net36),
    .A3(net132),
    .S0(net1021),
    .S1(clknet_1_1__leaf_net728),
    .X(net369));
 sky130_fd_sc_hd__mux4_1 c554 (.A0(net38),
    .A1(net154),
    .A2(net235),
    .A3(net947),
    .S0(clknet_1_1__leaf_net259),
    .S1(net984),
    .X(net370));
 sky130_fd_sc_hd__mux4_2 c555 (.A0(net359),
    .A1(net144),
    .A2(net264),
    .A3(net247),
    .S0(net244),
    .S1(net984),
    .X(net371));
 sky130_fd_sc_hd__mux4_1 c556 (.A0(net136),
    .A1(net358),
    .A2(net141),
    .A3(net580),
    .S0(net591),
    .S1(clknet_1_1__leaf_net726),
    .X(net372));
 sky130_fd_sc_hd__mux4_2 c557 (.A0(net792),
    .A1(net38),
    .A2(net120),
    .A3(net984),
    .S0(net800),
    .S1(net347),
    .X(net373));
 sky130_fd_sc_hd__mux4_1 c558 (.A0(net373),
    .A1(net792),
    .A2(net119),
    .A3(net1029),
    .S0(net665),
    .S1(net733),
    .X(net374));
 sky130_fd_sc_hd__mux4_1 c559 (.A0(net373),
    .A1(net348),
    .A2(net140),
    .A3(net568),
    .S0(net569),
    .S1(net594),
    .X(net375));
 sky130_fd_sc_hd__mux4_1 c560 (.A0(net355),
    .A1(net984),
    .A2(clknet_1_1__leaf_net368),
    .A3(net1012),
    .S0(clknet_1_1__leaf_net726),
    .S1(net735),
    .X(net376));
 sky130_fd_sc_hd__mux4_1 c561 (.A0(net960),
    .A1(net154),
    .A2(net1029),
    .A3(net246),
    .S0(net357),
    .S1(net735),
    .X(net377));
 sky130_fd_sc_hd__mux4_1 c562 (.A0(net377),
    .A1(net342),
    .A2(clknet_1_1__leaf_net376),
    .A3(net569),
    .S0(net591),
    .S1(net724),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 c563 (.A0(clknet_1_0__leaf_net361),
    .A1(net984),
    .A2(net377),
    .A3(net599),
    .S0(net990),
    .S1(net735),
    .X(net379));
 sky130_fd_sc_hd__mux4_1 c564 (.A0(net373),
    .A1(net377),
    .A2(net591),
    .A3(net729),
    .S0(net734),
    .S1(net736),
    .X(net380));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net1047),
    .A1(net984),
    .A2(net377),
    .A3(clknet_1_1__leaf_net728),
    .S0(net736),
    .S1(net737),
    .X(net381));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(clknet_1_1__leaf_net364),
    .A1(net661),
    .A2(net991),
    .A3(clknet_1_0__leaf_net875),
    .S0(net736),
    .S1(net737),
    .X(net382));
 sky130_fd_sc_hd__mux4_1 c567 (.A0(net1037),
    .A1(net614),
    .A2(clknet_1_1__leaf_net709),
    .A3(clknet_1_0__leaf_net875),
    .S0(net735),
    .S1(net737),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 c568 (.A0(net232),
    .A1(net272),
    .A2(clknet_1_1__leaf_net382),
    .A3(net984),
    .S0(net357),
    .S1(net735),
    .X(net384));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(net119),
    .A1(net357),
    .A2(net155),
    .A3(clknet_1_1__leaf_net384),
    .S0(net599),
    .S1(net733),
    .X(net385));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(clknet_1_1__leaf_net384),
    .A1(clknet_1_1__leaf_net383),
    .A3(net735),
    .S0(net737),
    .S1(net738),
    .X(net386));
 sky130_fd_sc_hd__mux4_1 c571 (.A0(net357),
    .A1(net614),
    .A2(clknet_1_1__leaf_net875),
    .A3(clknet_1_0__leaf_net728),
    .S0(net733),
    .S1(net738),
    .X(net387));
 sky130_fd_sc_hd__mux4_1 c572 (.A0(net889),
    .A1(net154),
    .A2(net1045),
    .A3(net808),
    .S0(net661),
    .S1(net688),
    .X(net388));
 sky130_fd_sc_hd__mux4_1 c573 (.A0(net154),
    .A1(net997),
    .A2(net824),
    .A3(net1003),
    .S0(net990),
    .S1(clknet_1_1__leaf_net690),
    .X(net880));
 sky130_fd_sc_hd__mux4_1 c574 (.A0(net286),
    .A1(net373),
    .A2(net71),
    .A3(net1008),
    .S0(net725),
    .S1(clknet_1_0__leaf_net726),
    .X(net389));
 sky130_fd_sc_hd__mux4_1 c575 (.A0(net808),
    .A1(clknet_1_0__leaf_net384),
    .A2(clknet_1_0__leaf_net300),
    .A3(net967),
    .S0(clknet_1_0__leaf_net287),
    .S1(net710),
    .X(net390));
 sky130_fd_sc_hd__mux4_1 c576 (.A0(clknet_1_1__leaf_net300),
    .A1(net1021),
    .A2(net803),
    .A3(net643),
    .S0(clknet_1_1__leaf_net689),
    .S1(net717),
    .X(net391));
 sky130_fd_sc_hd__mux4_2 c577 (.A0(net819),
    .A1(net569),
    .A2(net643),
    .A3(net718),
    .S0(net725),
    .S1(net730),
    .X(net890));
 sky130_fd_sc_hd__mux4_1 c578 (.A0(clknet_1_0__leaf_net384),
    .A1(net960),
    .A2(net824),
    .A3(net664),
    .S0(net992),
    .S1(net990),
    .X(net392));
 sky130_fd_sc_hd__mux4_2 c579 (.A0(net272),
    .A1(net1014),
    .A2(net1053),
    .A3(net243),
    .S0(net653),
    .S1(net725),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 c580 (.A0(clknet_1_1__leaf_net275),
    .A1(net1005),
    .A2(clknet_1_0__leaf_net383),
    .A3(clknet_1_1__leaf_net690),
    .S0(clknet_1_0__leaf_net728),
    .S1(net735),
    .X(net394));
 sky130_fd_sc_hd__mux4_1 c581 (.A0(net247),
    .A1(net288),
    .A2(net1003),
    .A3(net663),
    .S0(net992),
    .S1(net738),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(net979),
    .A1(net653),
    .A2(net658),
    .A3(net663),
    .S0(clknet_1_1__leaf_net690),
    .S1(clknet_1_0__leaf_net726),
    .X(net396));
 sky130_fd_sc_hd__mux4_1 c583 (.A0(clknet_1_1__leaf_net287),
    .A1(clknet_1_0__leaf_net396),
    .A2(net1014),
    .A3(net63),
    .S0(net568),
    .S1(net740),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 c584 (.A0(clknet_1_1__leaf_net382),
    .A1(net979),
    .A2(net247),
    .A3(net643),
    .S0(net718),
    .S1(clknet_1_0__leaf_net726),
    .X(net398));
 sky130_fd_sc_hd__mux4_1 c585 (.A0(net797),
    .A1(net824),
    .A2(net169),
    .A3(net884),
    .S0(net1009),
    .S1(net569),
    .X(net399));
 sky130_fd_sc_hd__mux4_1 c586 (.A0(net243),
    .A1(net234),
    .A2(clknet_1_0__leaf_net396),
    .A3(clknet_1_0__leaf_net728),
    .S0(net739),
    .S1(net743),
    .X(net887));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(net961),
    .A1(clknet_1_1__leaf_net398),
    .A2(clknet_1_1__leaf_net275),
    .A3(clknet_1_0__leaf_net259),
    .S0(net143),
    .S1(net658),
    .X(net400));
 sky130_fd_sc_hd__mux4_1 c588 (.A0(net357),
    .A1(net349),
    .A2(net947),
    .A3(net946),
    .S0(net731),
    .S1(net1078),
    .X(net401));
 sky130_fd_sc_hd__mux4_1 c589 (.A0(net36),
    .A1(clknet_1_0__leaf_net293),
    .A2(clknet_1_0__leaf_net880),
    .A3(clknet_1_0__leaf_net887),
    .S0(net614),
    .S1(net663),
    .X(net402));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(net136),
    .A1(net393),
    .A2(clknet_1_0__leaf_net887),
    .A3(clknet_1_0__leaf_net396),
    .S0(net974),
    .S1(clknet_1_0__leaf_net726),
    .X(net403));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(clknet_1_0__leaf_net383),
    .A1(net373),
    .A2(clknet_1_0__leaf_net396),
    .A3(net599),
    .S0(net719),
    .S1(net740),
    .X(net404));
 sky130_fd_sc_hd__sdfbbp_1 c592 (.CLK(clknet_4_9_0_clk),
    .D(clknet_1_1__leaf_net287),
    .RESET_B(net246),
    .SCD(net599),
    .SCE(net643),
    .SET_B(net1079),
    .Q(net406),
    .Q_N(net405));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(clknet_1_0__leaf_net887),
    .A1(net405),
    .A2(net797),
    .A3(net640),
    .S0(net643),
    .S1(net744),
    .X(net876));
 sky130_fd_sc_hd__mux4_1 c594 (.A0(clknet_1_0__leaf_net376),
    .A1(net60),
    .A2(net889),
    .A3(net393),
    .S0(net881),
    .S1(net696),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 c595 (.A0(net947),
    .A1(net54),
    .A2(clknet_1_0__leaf_net398),
    .A3(net846),
    .S0(net968),
    .S1(net722),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c596 (.A0(clknet_1_0__leaf_net277),
    .A1(net71),
    .A2(net1103),
    .A3(clknet_1_0__leaf_net306),
    .S0(net713),
    .S1(net720),
    .X(net409));
 sky130_fd_sc_hd__mux4_1 c597 (.A0(clknet_1_1__leaf_net185),
    .A1(net954),
    .A2(net888),
    .A3(net814),
    .S0(net646),
    .S1(net739),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 c598 (.A0(net408),
    .A1(net349),
    .A2(net888),
    .A3(net1024),
    .S0(net819),
    .S1(net736),
    .X(net411));
 sky130_fd_sc_hd__mux4_1 c599 (.A0(net371),
    .A1(net1029),
    .A2(net230),
    .A3(net948),
    .S0(net721),
    .S1(clknet_1_0__leaf_net746),
    .X(net412));
 sky130_fd_sc_hd__mux4_1 c600 (.A0(net970),
    .A1(net888),
    .A2(net846),
    .A3(net264),
    .S0(net723),
    .S1(net745),
    .X(net413));
 sky130_fd_sc_hd__mux4_2 c601 (.A0(clknet_1_0__leaf_net398),
    .A1(net974),
    .A2(clknet_1_1__leaf_net316),
    .A3(net1009),
    .S0(net143),
    .S1(net838),
    .X(net414));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(net412),
    .A1(net231),
    .A2(net406),
    .A3(net888),
    .S0(net838),
    .S1(clknet_1_0__leaf_net727),
    .X(net415));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(net890),
    .A1(net35),
    .A2(net60),
    .A3(net669),
    .S0(net988),
    .S1(clknet_1_0__leaf_net746),
    .X(net416));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(net890),
    .A1(net846),
    .A2(net1005),
    .A3(net936),
    .S0(net626),
    .S1(net646),
    .X(net417));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net270),
    .A1(net264),
    .A2(net231),
    .A3(net639),
    .S0(net669),
    .S1(net740),
    .X(net418));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net144),
    .A1(net61),
    .A2(clknet_1_0__leaf_net909),
    .A3(net1041),
    .S0(net120),
    .S1(net1011),
    .X(net419));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(clknet_1_0__leaf_net316),
    .A1(clknet_1_1__leaf_net416),
    .A2(net1085),
    .A3(net621),
    .S0(clknet_1_0__leaf_net727),
    .S1(net744),
    .X(net420));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net349),
    .A1(clknet_1_1__leaf_net278),
    .A2(net584),
    .A3(net624),
    .S0(net651),
    .S1(net736),
    .X(net421));
 sky130_fd_sc_hd__mux4_1 c609 (.A0(net417),
    .A1(net797),
    .A2(net936),
    .A3(net739),
    .S0(net745),
    .S1(clknet_1_0__leaf_net891),
    .X(net422));
 sky130_fd_sc_hd__mux4_1 c610 (.A0(net387),
    .A1(net58),
    .A2(net1051),
    .A3(net989),
    .S0(clknet_1_1__leaf_net746),
    .S1(clknet_1_0__leaf_net891),
    .X(net878));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net846),
    .A1(net624),
    .A2(clknet_1_0__leaf_net875),
    .A3(net711),
    .S0(net745),
    .S1(clknet_1_0__leaf_net891),
    .X(net423));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(clknet_1_0__leaf_net422),
    .A1(net418),
    .A2(net417),
    .A3(net803),
    .S0(net230),
    .S1(net651),
    .X(net424));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(clknet_1_0__leaf_net423),
    .A1(net1041),
    .A2(clknet_1_1__leaf_net422),
    .A3(net1024),
    .S0(net651),
    .S1(clknet_1_1__leaf_net746),
    .X(net425));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(clknet_1_1__leaf_net307),
    .A1(clknet_1_0__leaf_net878),
    .A2(net142),
    .A3(net639),
    .S0(clknet_1_0__leaf_net727),
    .S1(clknet_1_0__leaf_net891),
    .X(net426));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net425),
    .A1(net953),
    .A2(clknet_1_1__leaf_net423),
    .A3(net1027),
    .S0(net613),
    .S1(net745),
    .X(net427));
 sky130_fd_sc_hd__mux4_1 c616 (.A0(clknet_1_0__leaf_net416),
    .A1(net244),
    .A2(net918),
    .A3(net1012),
    .S0(net846),
    .S1(net702),
    .X(net428));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(net1045),
    .A1(clknet_1_0__leaf_net259),
    .A2(net985),
    .A3(net814),
    .S0(net801),
    .S1(clknet_1_1__leaf_net879),
    .X(net429));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(net71),
    .A1(clknet_1_0__leaf_net339),
    .A2(net58),
    .A3(net142),
    .S0(net858),
    .S1(net824),
    .X(net430));
 sky130_fd_sc_hd__mux4_1 c619 (.A0(net954),
    .A1(clknet_1_0__leaf_net325),
    .A2(net967),
    .A3(clknet_1_0__leaf_net382),
    .S0(net915),
    .S1(net747),
    .X(net431));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net797),
    .A1(net817),
    .A2(net1025),
    .A3(net919),
    .S0(net688),
    .S1(net893),
    .X(net873));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(net968),
    .A1(clknet_1_1__leaf_net339),
    .A2(net915),
    .A3(net625),
    .S0(net641),
    .S1(clknet_1_0__leaf_net891),
    .X(net432));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(net328),
    .A1(net819),
    .A2(net1016),
    .A3(net71),
    .S0(net667),
    .S1(net723),
    .X(net433));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(net888),
    .A1(net625),
    .A2(clknet_1_0__leaf_net649),
    .A3(net919),
    .S0(net893),
    .S1(net744),
    .X(net434));
 sky130_fd_sc_hd__mux4_1 c624 (.A0(net120),
    .A1(net824),
    .A2(net271),
    .A3(net888),
    .S0(net686),
    .S1(net1075),
    .X(net435));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net814),
    .A1(net433),
    .A2(clknet_1_1__leaf_net671),
    .A3(net744),
    .S0(clknet_1_0__leaf_net879),
    .S1(net749),
    .X(net436));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net296),
    .A1(net961),
    .A2(net1015),
    .A3(net1007),
    .S0(net1003),
    .S1(net989),
    .X(net437));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(clknet_1_0__leaf_net436),
    .A1(net405),
    .A2(net626),
    .A3(net638),
    .S0(net686),
    .S1(net866),
    .X(net438));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net393),
    .A1(net1025),
    .A2(net873),
    .A3(clknet_1_1__leaf_net330),
    .S0(clknet_1_0__leaf_net887),
    .S1(clknet_1_1__leaf_net649),
    .X(net439));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(net967),
    .A1(net968),
    .A2(net71),
    .A3(net296),
    .S0(clknet_1_1__leaf_net325),
    .S1(net702),
    .X(net440));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net440),
    .A1(net431),
    .A2(net846),
    .A3(net437),
    .S0(net747),
    .S1(net752),
    .X(net441));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(clknet_1_1__leaf_net338),
    .A1(net1027),
    .A2(clknet_1_1__leaf_net293),
    .A3(net1015),
    .S0(net657),
    .S1(clknet_1_0__leaf_net875),
    .X(net442));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net657),
    .A1(net677),
    .A2(net688),
    .A3(net700),
    .S0(net702),
    .S1(net752),
    .X(net867));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(net438),
    .A1(net437),
    .A2(net328),
    .A3(net657),
    .S0(net989),
    .S1(net751),
    .X(net443));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net406),
    .A1(net998),
    .A2(net433),
    .A3(net884),
    .S0(net437),
    .S1(net688),
    .X(net444));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net444),
    .A1(clknet_1_0__leaf_net325),
    .A2(net1087),
    .A3(clknet_1_0__leaf_net259),
    .S0(net1007),
    .S1(net919),
    .X(net445));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net803),
    .A1(net444),
    .A2(clknet_1_0__leaf_net339),
    .A3(net896),
    .S0(clknet_1_0__leaf_net649),
    .S1(net684),
    .X(net446));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net442),
    .A1(net443),
    .A2(clknet_1_0__leaf_net382),
    .A3(net633),
    .S0(clknet_1_1__leaf_net671),
    .S1(net700),
    .X(net447));
 sky130_fd_sc_hd__a41o_1 c660 (.A1(net777),
    .A2(net347),
    .A3(net1105),
    .A4(net996),
    .B1(net707),
    .X(net448));
 sky130_fd_sc_hd__mux4_1 c661 (.A0(clknet_1_1__leaf_net363),
    .A1(net997),
    .A2(net1033),
    .A3(net349),
    .S0(net951),
    .S1(net1023),
    .X(net449));
 sky130_fd_sc_hd__mux4_2 c662 (.A0(net241),
    .A1(net777),
    .A2(net964),
    .A3(net448),
    .S0(net127),
    .S1(net973),
    .X(net450));
 sky130_fd_sc_hd__a41o_1 c663 (.A1(net343),
    .A2(net342),
    .A3(net1003),
    .A4(net948),
    .B1(net707),
    .X(net451));
 sky130_fd_sc_hd__a41o_1 c664 (.A1(net1003),
    .A2(net996),
    .A3(net576),
    .A4(net642),
    .B1(net729),
    .X(net452));
 sky130_fd_sc_hd__a41o_1 c665 (.A1(net1057),
    .A2(net241),
    .A3(net568),
    .A4(net680),
    .B1(net684),
    .X(net453));
 sky130_fd_sc_hd__a41o_1 c666 (.A1(net450),
    .A2(net453),
    .A3(net965),
    .A4(net134),
    .B1(net981),
    .X(net454));
 sky130_fd_sc_hd__a41o_1 c667 (.A1(net128),
    .A2(net779),
    .A3(net454),
    .A4(net705),
    .B1(clknet_1_1__leaf_net727),
    .X(net455));
 sky130_fd_sc_hd__mux4_2 c668 (.A0(net134),
    .A1(net450),
    .A2(net1004),
    .A3(net965),
    .S0(net453),
    .S1(net654),
    .X(net456));
 sky130_fd_sc_hd__sdfbbn_1 c669 (.CLK_N(clknet_4_15_0_clk),
    .D(net242),
    .RESET_B(net342),
    .SCD(net456),
    .SCE(net568),
    .SET_B(net706),
    .Q(net458),
    .Q_N(net457));
 sky130_fd_sc_hd__mux4_1 c670 (.A0(net454),
    .A1(net965),
    .A2(net810),
    .A3(net127),
    .S0(net133),
    .S1(net654),
    .X(net459));
 sky130_fd_sc_hd__mux4_1 c671 (.A0(net1023),
    .A1(net1022),
    .A2(net457),
    .A3(net577),
    .S0(net704),
    .S1(net707),
    .X(net460));
 sky130_fd_sc_hd__sdfbbn_2 c672 (.CLK_N(clknet_4_15_0_clk),
    .D(net456),
    .RESET_B(net460),
    .SCD(net127),
    .SCE(net1023),
    .SET_B(net1074),
    .Q(net462),
    .Q_N(net461));
 sky130_fd_sc_hd__a41o_1 c673 (.A1(net346),
    .A2(net462),
    .A3(net456),
    .A4(net642),
    .B1(net1074),
    .X(net463));
 sky130_fd_sc_hd__a41o_2 c674 (.A1(net462),
    .A2(net981),
    .A3(net133),
    .A4(net1009),
    .B1(net655),
    .X(net464));
 sky130_fd_sc_hd__mux4_1 c675 (.A0(net453),
    .A1(net965),
    .A2(net462),
    .A3(net454),
    .S0(net464),
    .S1(net779),
    .X(net465));
 sky130_fd_sc_hd__mux4_1 c676 (.A0(net353),
    .A1(net448),
    .A2(net1014),
    .A3(net655),
    .S0(clknet_1_1__leaf_net727),
    .S1(net753),
    .X(net466));
 sky130_fd_sc_hd__mux4_1 c677 (.A0(net460),
    .A1(net464),
    .A2(net456),
    .A3(net461),
    .S0(clknet_1_1__leaf_net466),
    .S1(net958),
    .X(net467));
 sky130_fd_sc_hd__sdfbbp_1 c678 (.CLK(clknet_4_15_0_clk),
    .D(net448),
    .RESET_B(net464),
    .SCD(net456),
    .SCE(net991),
    .SET_B(net755),
    .Q(net469),
    .Q_N(net468));
 sky130_fd_sc_hd__mux4_1 c679 (.A0(net951),
    .A1(net468),
    .A2(net464),
    .A3(net454),
    .S1(net755),
    .X(net470));
 sky130_fd_sc_hd__mux4_2 c680 (.A0(net468),
    .A1(net464),
    .A2(net568),
    .A3(net577),
    .S0(net655),
    .S1(net755),
    .X(net471));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(net469),
    .A1(net461),
    .A2(net464),
    .A3(net450),
    .S0(net753),
    .S1(net755),
    .X(net472));
 sky130_fd_sc_hd__mux4_1 c682 (.A0(clknet_1_1__leaf_net365),
    .A1(net235),
    .A2(net1033),
    .A3(net456),
    .S0(net1032),
    .S1(net654),
    .X(net473));
 sky130_fd_sc_hd__mux4_1 c683 (.A0(net1037),
    .A1(net791),
    .A2(net242),
    .A3(net984),
    .S0(net960),
    .S1(net681),
    .X(net474));
 sky130_fd_sc_hd__mux4_1 c684 (.A0(net155),
    .A1(net983),
    .A2(net1063),
    .A3(net619),
    .S0(net736),
    .S1(net754),
    .X(net475));
 sky130_fd_sc_hd__mux4_1 c685 (.A0(net348),
    .A1(net469),
    .A2(net464),
    .A3(net985),
    .S0(net42),
    .S1(net681),
    .X(net476));
 sky130_fd_sc_hd__mux4_1 c686 (.A0(net1023),
    .A1(net1026),
    .A2(clknet_1_1__leaf_net278),
    .A3(net1022),
    .S0(net245),
    .S1(net756),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c687 (.A0(net464),
    .A1(net469),
    .A2(net371),
    .A3(clknet_1_1__leaf_net709),
    .S0(net738),
    .S1(net757),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c688 (.A0(net1009),
    .A1(net779),
    .A2(net791),
    .A3(net155),
    .S0(net468),
    .S1(net771),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c689 (.A0(net469),
    .A1(net371),
    .A2(net1026),
    .A3(net464),
    .S0(net456),
    .S1(net1016),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c690 (.A0(net958),
    .A1(net134),
    .A2(clknet_1_0__leaf_net466),
    .A3(net946),
    .S0(net971),
    .S1(net630),
    .X(net481));
 sky130_fd_sc_hd__mux4_1 c691 (.A0(net1023),
    .A1(net1006),
    .A2(net619),
    .A3(net724),
    .S0(net729),
    .S1(net758),
    .X(net482));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(net39),
    .A1(net766),
    .A2(clknet_1_1__leaf_net278),
    .A3(net452),
    .S0(net342),
    .S1(net754),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c693 (.A0(clknet_1_0__leaf_net466),
    .A1(net352),
    .A2(net371),
    .A3(net242),
    .S0(net779),
    .S1(net760),
    .X(net484));
 sky130_fd_sc_hd__mux4_1 c694 (.A0(net1004),
    .A1(net1022),
    .A2(net1025),
    .A3(net630),
    .S0(net642),
    .S1(net758),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c695 (.A0(net456),
    .A1(net1032),
    .A2(net636),
    .A3(net734),
    .S0(net759),
    .S1(net760),
    .X(net486));
 sky130_fd_sc_hd__mux4_1 c696 (.A0(net482),
    .A1(net791),
    .A2(clknet_1_1__leaf_net709),
    .A3(net732),
    .S0(net754),
    .S1(net760),
    .X(net487));
 sky130_fd_sc_hd__mux4_1 c697 (.A0(clknet_1_1__leaf_net484),
    .A1(clknet_1_1__leaf_net364),
    .A2(net1032),
    .A3(net983),
    .S0(net754),
    .S1(net761),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(net487),
    .A1(net461),
    .A2(net468),
    .A3(net730),
    .S0(net756),
    .S1(net760),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(net157),
    .A1(net983),
    .A2(net580),
    .A3(net661),
    .S0(net705),
    .S1(net734),
    .X(net490));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net155),
    .A1(net47),
    .A2(net234),
    .A3(net926),
    .S0(net759),
    .S1(net761),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(net456),
    .A1(net469),
    .A2(clknet_1_0__leaf_net484),
    .A3(clknet_1_1__leaf_net478),
    .S0(net631),
    .S1(net753),
    .X(net492));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net464),
    .A1(net342),
    .A2(net799),
    .A3(net1016),
    .S0(net631),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(net474),
    .A1(net157),
    .A2(net1026),
    .A3(net985),
    .S0(net636),
    .S1(net926),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net476),
    .A1(net1033),
    .A2(net245),
    .A3(net1022),
    .S0(net730),
    .S1(net740),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(clknet_1_0__leaf_net365),
    .A1(net39),
    .A2(net458),
    .A3(clknet_1_1__leaf_net396),
    .S0(net643),
    .S1(net738),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c706 (.A0(net472),
    .A1(net1025),
    .A2(net40),
    .A3(net817),
    .S0(net782),
    .S1(net805),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c707 (.A0(net802),
    .A1(net169),
    .A2(net632),
    .A3(clknet_1_1__leaf_net689),
    .S0(net711),
    .S1(net741),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(clknet_1_0__leaf_net396),
    .A1(clknet_1_1__leaf_net293),
    .A2(net652),
    .A3(net705),
    .S0(net743),
    .S1(net762),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(net462),
    .A1(net791),
    .A2(net802),
    .A3(clknet_1_1__leaf_net499),
    .S0(clknet_1_1__leaf_net489),
    .S1(net760),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net452),
    .A1(net800),
    .A2(clknet_1_1__leaf_net689),
    .A3(net705),
    .S0(net718),
    .S1(net736),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net802),
    .A1(clknet_1_0__leaf_net396),
    .A2(net34),
    .A3(net981),
    .S0(net666),
    .S1(net762),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net286),
    .A1(clknet_1_0__leaf_net489),
    .A2(net472),
    .A3(clknet_1_1__leaf_net293),
    .S0(net39),
    .S1(net753),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c713 (.A0(net974),
    .A1(net984),
    .A2(net640),
    .A3(net663),
    .S0(net724),
    .S1(net763),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(net157),
    .A1(net342),
    .A2(net805),
    .A3(net462),
    .S0(net264),
    .S1(net680),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net458),
    .A1(clknet_1_1__leaf_net396),
    .A2(net765),
    .A3(net744),
    .S0(net762),
    .S1(net763),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net802),
    .A1(net985),
    .A2(net342),
    .A3(net457),
    .S0(net992),
    .S1(net874),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net1065),
    .A1(net817),
    .A2(net256),
    .A3(clknet_1_0__leaf_net499),
    .S0(net271),
    .S1(net647),
    .X(net508));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(clknet_1_1__leaf_net506),
    .A1(net663),
    .A2(net736),
    .A3(net753),
    .S0(net757),
    .S1(net762),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(clknet_1_1__leaf_net396),
    .A1(net448),
    .A2(clknet_1_0__leaf_net506),
    .A3(net1022),
    .S0(net771),
    .S1(clknet_1_1__leaf_net709),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net500),
    .A1(net504),
    .A2(clknet_1_0__leaf_net506),
    .A3(net981),
    .S0(net663),
    .S1(net874),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net511),
    .A1(net777),
    .A2(clknet_1_0__leaf_net365),
    .A3(clknet_1_1__leaf_net499),
    .S0(net774),
    .S1(net1007),
    .X(net512));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(clknet_1_0__leaf_net478),
    .A1(net510),
    .A2(clknet_1_1__leaf_net496),
    .A3(net946),
    .S0(net774),
    .S1(net717),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net256),
    .A1(clknet_1_1__leaf_net496),
    .A2(clknet_1_1__leaf_net506),
    .A3(net461),
    .S0(net983),
    .S1(net762),
    .X(net514));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(clknet_1_0__leaf_net496),
    .A1(net642),
    .A2(net652),
    .A3(net658),
    .S0(net680),
    .S1(net763),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net169),
    .A1(net371),
    .A2(net633),
    .A3(net652),
    .S0(clknet_1_0__leaf_net691),
    .S1(net763),
    .X(net516));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net846),
    .A1(net965),
    .A2(net642),
    .A3(net705),
    .S0(net711),
    .S1(net738),
    .X(net517));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net197),
    .A1(net800),
    .A2(net926),
    .A3(net989),
    .S0(clknet_1_0__leaf_net727),
    .S1(clknet_1_0__leaf_net764),
    .X(net518));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net965),
    .A1(net958),
    .A2(net245),
    .A3(clknet_1_1__leaf_net691),
    .S0(net731),
    .S1(net741),
    .X(net519));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(net485),
    .A1(net948),
    .A2(net952),
    .A3(net1011),
    .S0(net641),
    .S1(net642),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net805),
    .A1(clknet_1_1__leaf_net306),
    .A2(net245),
    .A3(net661),
    .S0(net684),
    .S1(clknet_1_0__leaf_net727),
    .X(net521));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(clknet_1_0__leaf_net496),
    .A1(net838),
    .A2(net600),
    .A3(net648),
    .S0(clknet_1_1__leaf_net671),
    .S1(net763),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(clknet_1_1__leaf_net278),
    .A1(clknet_1_0__leaf_net427),
    .A2(clknet_1_0__leaf_net496),
    .A3(clknet_1_0__leaf_net868),
    .S0(clknet_1_1__leaf_net306),
    .S1(net989),
    .X(net523));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net765),
    .A1(net190),
    .A2(net838),
    .A3(clknet_1_0__leaf_net424),
    .S0(net800),
    .S1(net42),
    .X(net524));
 sky130_fd_sc_hd__mux4_2 c734 (.A0(net791),
    .A1(net40),
    .A2(net980),
    .A3(clknet_1_1__leaf_net650),
    .S0(net661),
    .S1(net763),
    .X(net525));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net63),
    .A1(net632),
    .A2(clknet_1_1__leaf_net650),
    .A3(net738),
    .S0(net756),
    .S1(clknet_1_1__leaf_net764),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(net1025),
    .A1(net838),
    .A2(clknet_1_1__leaf_net526),
    .A3(net577),
    .S0(clknet_1_0__leaf_net727),
    .S1(net761),
    .X(net527));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net520),
    .A1(net471),
    .A2(net877),
    .A3(net681),
    .S0(net732),
    .S1(clknet_1_1__leaf_net764),
    .X(net528));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net83),
    .A1(net235),
    .A2(clknet_1_1__leaf_net304),
    .A3(net633),
    .S0(net741),
    .S1(net762),
    .X(net529));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(net482),
    .A1(net520),
    .A2(net245),
    .A3(net624),
    .S0(net681),
    .S1(net684),
    .X(net530));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(net524),
    .A1(clknet_1_0__leaf_net526),
    .A2(net319),
    .A3(clknet_1_1__leaf_net427),
    .S0(net765),
    .S1(clknet_1_1__leaf_net891),
    .X(net531));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(net509),
    .A1(net765),
    .A2(net971),
    .A3(net926),
    .S0(net665),
    .S1(net989),
    .X(net532));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(clknet_1_0__leaf_net532),
    .A1(clknet_1_0__leaf_net499),
    .A2(net838),
    .A3(net870),
    .S0(clknet_1_1__leaf_net691),
    .S1(net757),
    .X(net533));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(net485),
    .A1(net872),
    .A2(clknet_1_1__leaf_net532),
    .A3(net958),
    .S0(net600),
    .S1(net870),
    .X(net534));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(net471),
    .A1(clknet_1_1__leaf_net527),
    .A2(clknet_1_1__leaf_net532),
    .A3(net985),
    .S0(net661),
    .S1(net763),
    .X(net535));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(net47),
    .A1(clknet_1_0__leaf_net532),
    .A2(net645),
    .A3(clknet_1_0__leaf_net727),
    .S0(net741),
    .S1(clknet_1_0__leaf_net764),
    .X(net536));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(clknet_1_1__leaf_net304),
    .A1(clknet_1_1__leaf_net424),
    .A2(net536),
    .A3(clknet_1_0__leaf_net527),
    .S0(clknet_1_0__leaf_net532),
    .S1(net870),
    .X(net537));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(clknet_1_1__leaf_net304),
    .A1(net983),
    .A2(net632),
    .A3(net648),
    .S0(net991),
    .S1(net763),
    .X(net538));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net796),
    .A1(net433),
    .A2(net518),
    .A3(net985),
    .S0(net54),
    .S1(net656),
    .X(net539));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net1007),
    .A1(net1003),
    .A2(net858),
    .A3(net613),
    .S0(net637),
    .S1(net656),
    .X(net540));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(clknet_1_0__leaf_net364),
    .A1(net43),
    .A2(net1085),
    .A3(clknet_1_1__leaf_net649),
    .S0(clknet_1_0__leaf_net650),
    .S1(net667),
    .X(net541));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(clknet_1_0__leaf_net382),
    .A1(net235),
    .A2(net805),
    .A3(net799),
    .S0(net1011),
    .S1(clknet_1_1__leaf_net689),
    .X(net542));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net538),
    .A1(net952),
    .A2(clknet_1_1__leaf_net436),
    .A3(net633),
    .S0(net637),
    .S1(net665),
    .X(net543));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net540),
    .A1(clknet_1_0__leaf_net364),
    .A2(net817),
    .A3(clknet_1_1__leaf_net649),
    .S0(net684),
    .S1(net736),
    .X(net544));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net264),
    .A1(net981),
    .A2(clknet_1_1__leaf_net525),
    .A3(net638),
    .S0(clknet_1_0__leaf_net650),
    .S1(net762),
    .X(net545));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net1064),
    .A1(clknet_1_1__leaf_net293),
    .A2(net1022),
    .A3(net774),
    .S0(net988),
    .S1(net756),
    .X(net546));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net54),
    .A1(clknet_1_0__leaf_net525),
    .A2(net774),
    .A3(net858),
    .S0(net989),
    .S1(net866),
    .X(net547));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net501),
    .A1(net42),
    .A2(clknet_1_0__leaf_net547),
    .A3(net953),
    .S0(net789),
    .S1(net762),
    .X(net548));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(clknet_1_1__leaf_net306),
    .A1(net800),
    .A2(net545),
    .A3(net29),
    .S0(net624),
    .S1(net665),
    .X(net549));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net805),
    .A1(net544),
    .A2(net771),
    .A3(clknet_1_1__leaf_net691),
    .S0(net745),
    .S1(net748),
    .X(net550));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net502),
    .A1(net771),
    .A2(net29),
    .A3(net546),
    .S0(clknet_1_1__leaf_net689),
    .S1(net748),
    .X(net551));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net948),
    .A1(net1009),
    .A2(net551),
    .A3(clknet_1_1__leaf_net529),
    .S0(net1066),
    .S1(net631),
    .X(net552));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net953),
    .A1(net1011),
    .A2(net543),
    .A3(net43),
    .S0(net645),
    .S1(net744),
    .X(net553));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(net319),
    .A1(net1044),
    .A2(net552),
    .A3(net1003),
    .S0(net656),
    .S1(net717),
    .X(net554));
 sky130_fd_sc_hd__mux4_1 c764 (.A0(net349),
    .A1(net1012),
    .A2(clknet_1_1__leaf_net691),
    .A3(net988),
    .S0(net745),
    .S1(net757),
    .X(net555));
 sky130_fd_sc_hd__mux4_1 c765 (.A0(net245),
    .A1(clknet_1_1__leaf_net547),
    .A2(net629),
    .A3(net648),
    .S0(clknet_1_1__leaf_net671),
    .S1(net761),
    .X(net556));
 sky130_fd_sc_hd__a41o_1 c766 (.A1(net846),
    .A2(clknet_1_0__leaf_net529),
    .A3(net539),
    .A4(net926),
    .B1(net667),
    .X(net557));
 sky130_fd_sc_hd__mux4_1 c767 (.A0(net542),
    .A1(net550),
    .A2(net641),
    .A3(net645),
    .S0(net700),
    .S1(net761),
    .X(net558));
 sky130_fd_sc_hd__mux4_1 c768 (.A0(net799),
    .A1(net533),
    .A2(net558),
    .A3(net629),
    .S0(net645),
    .S1(net750),
    .X(net559));
 sky130_fd_sc_hd__mux4_1 c769 (.A0(net271),
    .A1(net517),
    .A2(net34),
    .A3(net559),
    .S0(net877),
    .S1(net631),
    .X(net560));
 sky130_fd_sc_hd__xnor2_1 merge790 (.A(net429),
    .B(net439),
    .Y(net561));
 sky130_fd_sc_hd__xnor2_1 merge791 (.A(net481),
    .B(net486),
    .Y(net562));
 sky130_fd_sc_hd__xnor2_1 merge792 (.A(net208),
    .B(net189),
    .Y(net563));
 sky130_fd_sc_hd__dfrbp_2 merge793 (.CLK(clknet_4_1_0_clk),
    .D(net86),
    .RESET_B(net90),
    .Q(net898),
    .Q_N(net564));
 sky130_fd_sc_hd__dfrbp_2 merge794 (.CLK(clknet_4_5_0_clk),
    .D(net44),
    .Q(net49),
    .Q_N(net565));
 sky130_fd_sc_hd__xnor2_1 merge795 (.A(net519),
    .B(net521),
    .Y(net567));
 sky130_fd_sc_hd__dfrtn_1 merge796 (.CLK_N(clknet_4_13_0_clk),
    .D(net350),
    .RESET_B(net344),
    .Q(net568));
 sky130_fd_sc_hd__dfrtp_2 merge797 (.CLK(clknet_4_12_0_clk),
    .D(net369),
    .RESET_B(net370),
    .Q(net569));
 sky130_fd_sc_hd__xnor2_1 merge798 (.A(net324),
    .B(net326),
    .Y(net570));
 sky130_fd_sc_hd__xnor2_2 merge799 (.A(net409),
    .B(net414),
    .Y(net571));
 sky130_fd_sc_hd__xnor2_1 merge800 (.A(net170),
    .B(net173),
    .Y(net572));
 sky130_fd_sc_hd__dfrtp_4 merge801 (.CLK(clknet_4_6_0_clk),
    .D(net156),
    .RESET_B(net164),
    .Q(net573));
 sky130_fd_sc_hd__dfrtp_1 merge802 (.CLK(clknet_4_3_0_clk),
    .D(net305),
    .RESET_B(net309),
    .Q(net574));
 sky130_fd_sc_hd__xnor2_1 merge803 (.A(net209),
    .B(net217),
    .Y(net575));
 sky130_fd_sc_hd__dfsbp_1 merge804 (.CLK(clknet_4_15_0_clk),
    .SET_B(net449),
    .Q(net577),
    .Q_N(net470));
 sky130_fd_sc_hd__dfsbp_2 merge805 (.CLK(clknet_4_1_0_clk),
    .D(net65),
    .Q(net72),
    .Q_N(net578));
 sky130_fd_sc_hd__dfstp_1 merge806 (.CLK(clknet_4_0_0_clk),
    .D(net115),
    .SET_B(net114),
    .Q(net933));
 sky130_fd_sc_hd__dfstp_2 merge807 (.CLK(clknet_4_6_0_clk),
    .D(net279),
    .SET_B(net266),
    .Q(net580));
 sky130_fd_sc_hd__xnor2_1 merge808 (.A(net497),
    .B(net498),
    .Y(net581));
 sky130_fd_sc_hd__dfstp_2 merge809 (.CLK(clknet_4_7_0_clk),
    .D(net233),
    .SET_B(net249),
    .Q(net582));
 sky130_fd_sc_hd__dlrbn_2 merge810 (.D(net138),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net125),
    .Q(net584),
    .Q_N(net583));
 sky130_fd_sc_hd__xnor2_1 merge811 (.A(net111),
    .B(net112),
    .Y(net585));
 sky130_fd_sc_hd__xnor2_1 merge812 (.A(net560),
    .B(net541),
    .Y(net586));
 sky130_fd_sc_hd__xnor2_1 merge813 (.A(net285),
    .B(net298),
    .Y(net587));
 sky130_fd_sc_hd__xnor2_1 merge814 (.A(net391),
    .B(net395),
    .Y(net588));
 sky130_fd_sc_hd__xnor2_1 merge815 (.A(net492),
    .B(net490),
    .Y(net589));
 sky130_fd_sc_hd__dlrbn_2 merge816 (.D(net162),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net129),
    .Q(net591),
    .Q_N(net590));
 sky130_fd_sc_hd__dlrbp_2 merge817 (.D(net91),
    .GATE(clknet_4_1_0_clk),
    .Q(net92),
    .Q_N(net901));
 sky130_fd_sc_hd__xnor2_1 merge818 (.A(net488),
    .B(net378),
    .Y(net593));
 sky130_fd_sc_hd__dlrbp_2 merge819 (.D(net51),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net46),
    .Q(net877),
    .Q_N(net594));
 sky130_fd_sc_hd__xnor2_1 merge820 (.A(net227),
    .B(net225),
    .Y(net595));
 sky130_fd_sc_hd__xnor2_1 merge821 (.A(net175),
    .B(net188),
    .Y(net596));
 sky130_fd_sc_hd__xnor2_1 merge822 (.A(net415),
    .B(net447),
    .Y(net597));
 sky130_fd_sc_hd__dlrtn_2 merge823 (.D(net105),
    .GATE_N(clknet_4_0_0_clk),
    .RESET_B(net116),
    .Q(net915));
 sky130_fd_sc_hd__dlrtn_2 merge824 (.D(net101),
    .GATE_N(clknet_4_0_0_clk),
    .RESET_B(net585),
    .Q(net882));
 sky130_fd_sc_hd__dlrtn_1 merge825 (.D(net68),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net70));
 sky130_fd_sc_hd__dlrtp_1 merge826 (.D(net402),
    .GATE(clknet_4_12_0_clk),
    .RESET_B(net374),
    .Q(net599));
 sky130_fd_sc_hd__dlrtp_1 merge827 (.D(net66),
    .GATE(clknet_4_4_0_clk),
    .Q(net67));
 sky130_fd_sc_hd__xnor2_1 merge828 (.A(net595),
    .B(net445),
    .Y(net601));
 sky130_fd_sc_hd__xnor2_1 merge829 (.A(net221),
    .B(net219),
    .Y(net602));
 sky130_fd_sc_hd__xnor2_1 merge830 (.A(net340),
    .B(net333),
    .Y(net603));
 sky130_fd_sc_hd__xnor2_1 merge831 (.A(net426),
    .B(net537),
    .Y(net604));
 sky130_fd_sc_hd__xnor2_1 merge832 (.A(net586),
    .B(net557),
    .Y(net605));
 sky130_fd_sc_hd__xnor2_1 merge833 (.A(net331),
    .B(net329),
    .Y(net606));
 sky130_fd_sc_hd__xnor2_1 merge834 (.A(net421),
    .B(net556),
    .Y(net607));
 sky130_fd_sc_hd__xnor2_1 merge835 (.A(net548),
    .B(net549),
    .Y(net608));
 sky130_fd_sc_hd__dlrtp_1 merge836 (.D(net561),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net413),
    .Q(net936));
 sky130_fd_sc_hd__xnor2_1 merge837 (.A(net522),
    .B(net555),
    .Y(net609));
 sky130_fd_sc_hd__xnor2_1 merge838 (.A(net516),
    .B(net515),
    .Y(net610));
 sky130_fd_sc_hd__xnor2_1 merge839 (.A(net507),
    .B(net508),
    .Y(net611));
 sky130_fd_sc_hd__xnor2_1 merge840 (.A(net512),
    .B(net611),
    .Y(net612));
 sky130_fd_sc_hd__edfxbp_1 merge841 (.CLK(clknet_4_8_0_clk),
    .D(net315),
    .DE(net604),
    .Q(net897),
    .Q_N(net613));
 sky130_fd_sc_hd__edfxtp_1 merge842 (.CLK(clknet_4_14_0_clk),
    .DE(net381),
    .Q(net386));
 sky130_fd_sc_hd__sdlclkp_1 merge843 (.CLK(clknet_4_12_0_clk),
    .SCE(net280),
    .GCLK(net281));
 sky130_fd_sc_hd__sdlclkp_2 merge844 (.CLK(clknet_4_6_0_clk),
    .GATE(net186),
    .SCE(net596),
    .GCLK(net911));
 sky130_fd_sc_hd__xnor2_1 merge845 (.A(net553),
    .B(net554),
    .Y(net616));
 sky130_fd_sc_hd__sdlclkp_4 merge846 (.CLK(clknet_4_2_0_clk),
    .GATE(net323),
    .SCE(net603),
    .GCLK(net894));
 sky130_fd_sc_hd__xnor2_1 merge847 (.A(net216),
    .B(net226),
    .Y(net617));
 sky130_fd_sc_hd__dfrbp_2 merge848 (.CLK(clknet_4_9_0_clk),
    .D(net274),
    .RESET_B(net587),
    .Q(net619),
    .Q_N(net618));
 sky130_fd_sc_hd__xnor2_1 merge849 (.A(net535),
    .B(net534),
    .Y(net620));
 sky130_fd_sc_hd__dfrbp_1 merge850 (.CLK(clknet_4_3_0_clk),
    .D(net310),
    .RESET_B(net312),
    .Q(net622),
    .Q_N(net621));
 sky130_fd_sc_hd__xnor2_1 merge851 (.A(net616),
    .B(net567),
    .Y(net623));
 sky130_fd_sc_hd__dfrtn_1 merge852 (.CLK_N(clknet_4_2_0_clk),
    .D(net606),
    .RESET_B(net601),
    .Q(net896));
 sky130_fd_sc_hd__dfrtp_2 merge853 (.CLK(clknet_4_9_0_clk),
    .D(net407),
    .RESET_B(net597),
    .Q(net624));
 sky130_fd_sc_hd__dfrtp_1 merge854 (.CLK(clknet_4_2_0_clk),
    .D(net570),
    .RESET_B(net341),
    .Q(net625));
 sky130_fd_sc_hd__dfrtp_4 merge855 (.CLK(clknet_4_2_0_clk),
    .D(net193),
    .RESET_B(net321),
    .Q(net626));
 sky130_fd_sc_hd__dfsbp_1 merge856 (.CLK(clknet_4_0_0_clk),
    .D(net322),
    .SET_B(net602),
    .Q(net628),
    .Q_N(net627));
 sky130_fd_sc_hd__dfsbp_1 merge857 (.CLK(clknet_4_11_0_clk),
    .D(net480),
    .SET_B(net605),
    .Q(net630),
    .Q_N(net629));
 sky130_fd_sc_hd__dfstp_2 merge858 (.CLK(clknet_4_10_0_clk),
    .D(net491),
    .SET_B(net608),
    .Q(net631));
 sky130_fd_sc_hd__dfstp_1 merge859 (.CLK(clknet_4_14_0_clk),
    .SET_B(net589),
    .Q(net493));
 sky130_fd_sc_hd__dfstp_1 merge860 (.CLK(clknet_4_10_0_clk),
    .D(net610),
    .SET_B(net446),
    .Q(net633));
 sky130_fd_sc_hd__dlrbn_1 merge861 (.D(net575),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net198),
    .Q(net635),
    .Q_N(net634));
 sky130_fd_sc_hd__dlrbn_1 merge862 (.D(net581),
    .GATE_N(clknet_4_11_0_clk),
    .RESET_B(net562),
    .Q(net637),
    .Q_N(net636));
 sky130_fd_sc_hd__dlrbp_1 merge863 (.D(net571),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net435),
    .Q(net639),
    .Q_N(net638));
 sky130_fd_sc_hd__dlrbp_2 merge864 (.D(net607),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net400),
    .Q(net641),
    .Q_N(net640));
 sky130_fd_sc_hd__dlrtn_2 merge865 (.D(net451),
    .GATE_N(clknet_4_14_0_clk),
    .RESET_B(net612),
    .Q(net642));
 sky130_fd_sc_hd__dlrtn_2 merge866 (.D(net213),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net201),
    .Q(net902));
 sky130_fd_sc_hd__dlrtn_2 merge867 (.D(net388),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net404),
    .Q(net643));
 sky130_fd_sc_hd__dlrtp_2 merge868 (.D(net215),
    .GATE(clknet_4_0_0_clk),
    .RESET_B(net220),
    .Q(net644));
 sky130_fd_sc_hd__dlrtp_1 merge869 (.D(net620),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net609),
    .Q(net645));
 sky130_fd_sc_hd__dlrtp_2 merge870 (.D(net207),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net205),
    .Q(net646));
 sky130_fd_sc_hd__edfxbp_1 merge871 (.CLK(clknet_4_3_0_clk),
    .D(net302),
    .DE(net295),
    .Q(net648),
    .Q_N(net647));
 sky130_fd_sc_hd__edfxtp_1 merge872 (.CLK(clknet_4_10_0_clk),
    .D(net531),
    .DE(net530),
    .Q(net870));
 sky130_fd_sc_hd__sdlclkp_1 merge873 (.CLK(clknet_4_2_0_clk),
    .GATE(net229),
    .SCE(net223),
    .GCLK(net649));
 sky130_fd_sc_hd__sdlclkp_2 merge874 (.CLK(clknet_4_2_0_clk),
    .GATE(net617),
    .SCE(net200),
    .GCLK(net925));
 sky130_fd_sc_hd__sdlclkp_4 merge875 (.CLK(clknet_4_10_0_clk),
    .GATE(net528),
    .SCE(net523),
    .GCLK(net650));
 sky130_fd_sc_hd__dfrbp_1 merge876 (.CLK(clknet_4_11_0_clk),
    .D(net495),
    .RESET_B(net419),
    .Q(net652),
    .Q_N(net651));
 sky130_fd_sc_hd__dfrbp_2 merge877 (.CLK(clknet_4_13_0_clk),
    .D(net455),
    .RESET_B(net588),
    .Q(net654),
    .Q_N(net653));
 sky130_fd_sc_hd__dfrtn_1 merge878 (.CLK_N(clknet_4_10_0_clk),
    .D(net463),
    .RESET_B(net320),
    .Q(net655));
 sky130_fd_sc_hd__dfrtp_4 merge879 (.CLK(clknet_4_11_0_clk),
    .D(net623),
    .RESET_B(net477),
    .Q(net926));
 sky130_fd_sc_hd__dfrtp_4 merge880 (.CLK(clknet_4_8_0_clk),
    .D(net337),
    .RESET_B(net318),
    .Q(net656));
 sky130_fd_sc_hd__dfrtp_4 merge881 (.CLK(clknet_4_2_0_clk),
    .D(net336),
    .RESET_B(net563),
    .Q(net919));
 sky130_fd_sc_hd__dfsbp_2 merge882 (.CLK(clknet_4_8_0_clk),
    .D(net392),
    .SET_B(net441),
    .Q(net658),
    .Q_N(net657));
 sky130_fd_sc_hd__dfsbp_2 merge883 (.CLK(clknet_4_4_0_clk),
    .D(net572),
    .SET_B(net178),
    .Q(net660),
    .Q_N(net659));
 sky130_fd_sc_hd__dfstp_2 merge884 (.CLK(clknet_4_14_0_clk),
    .D(net513),
    .SET_B(net593),
    .Q(net661));
 sky130_fd_sc_hd__dfstp_2 merge885 (.CLK(clknet_4_2_0_clk),
    .D(net204),
    .SET_B(net228),
    .Q(net662));
 sky130_fd_sc_hd__dfstp_1 merge886 (.CLK(clknet_4_12_0_clk),
    .D(net403),
    .SET_B(net394),
    .Q(net663));
 sky130_fd_sc_hd__dfxbp_2 s887 (.CLK(clknet_4_4_0_clk),
    .D(net50),
    .Q(net665),
    .Q_N(net664));
 sky130_fd_sc_hd__dfxbp_2 s888 (.CLK(clknet_4_1_0_clk),
    .D(net69),
    .Q(net667),
    .Q_N(net666));
 sky130_fd_sc_hd__dfxtp_1 s889 (.CLK(clknet_4_1_0_clk),
    .D(net73),
    .Q(net668));
 sky130_fd_sc_hd__dfxtp_2 s890 (.CLK(clknet_4_1_0_clk),
    .D(net75),
    .Q(net669));
 sky130_fd_sc_hd__dfxtp_4 s891 (.CLK(clknet_4_1_0_clk),
    .D(net76),
    .Q(net670));
 sky130_fd_sc_hd__dlclkp_1 s892 (.CLK(clknet_4_1_0_clk),
    .GATE(net77),
    .GCLK(net671));
 sky130_fd_sc_hd__dlclkp_2 s893 (.CLK(clknet_4_1_0_clk),
    .GATE(net93),
    .GCLK(net672));
 sky130_fd_sc_hd__dlclkp_4 s894 (.CLK(clknet_4_0_0_clk),
    .GATE(net95),
    .GCLK(net673));
 sky130_fd_sc_hd__dlxbn_1 s895 (.D(net97),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net675),
    .Q_N(net674));
 sky130_fd_sc_hd__dlxbn_1 s896 (.D(net99),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net677),
    .Q_N(net676));
 sky130_fd_sc_hd__dlxbp_1 s897 (.D(net102),
    .GATE(clknet_4_0_0_clk),
    .Q(net885),
    .Q_N(net678));
 sky130_fd_sc_hd__dlxtn_2 s898 (.D(net106),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net679));
 sky130_fd_sc_hd__dlxtn_1 s899 (.D(net109),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net934));
 sky130_fd_sc_hd__dlxtn_2 s900 (.D(net126),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net680));
 sky130_fd_sc_hd__dlxtp_1 s901 (.D(net135),
    .GATE(clknet_4_7_0_clk),
    .Q(net681));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s902 (.D(net137),
    .SLEEP_B(clknet_4_7_0_clk),
    .Q(net682));
 sky130_fd_sc_hd__dfxbp_2 s903 (.CLK(clknet_4_7_0_clk),
    .D(net139),
    .Q(net684),
    .Q_N(net683));
 sky130_fd_sc_hd__dfxbp_2 s904 (.CLK(clknet_4_4_0_clk),
    .D(net151),
    .Q(net686),
    .Q_N(net685));
 sky130_fd_sc_hd__dfxtp_2 s905 (.CLK(clknet_4_5_0_clk),
    .D(net152),
    .Q(net687));
 sky130_fd_sc_hd__dfxtp_4 s906 (.CLK(clknet_4_5_0_clk),
    .D(net159),
    .Q(net688));
 sky130_fd_sc_hd__dfxtp_2 s907 (.CLK(clknet_4_4_0_clk),
    .D(net172),
    .Q(net899));
 sky130_fd_sc_hd__dlclkp_1 s908 (.CLK(clknet_4_4_0_clk),
    .GATE(net177),
    .GCLK(net689));
 sky130_fd_sc_hd__dlclkp_2 s909 (.CLK(clknet_4_1_0_clk),
    .GATE(net179),
    .GCLK(net690));
 sky130_fd_sc_hd__dlclkp_4 s910 (.CLK(clknet_4_6_0_clk),
    .GATE(net180),
    .GCLK(net691));
 sky130_fd_sc_hd__dlxbn_1 s911 (.D(net181),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net693),
    .Q_N(net692));
 sky130_fd_sc_hd__dlxbn_1 s912 (.D(net182),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net695),
    .Q_N(net694));
 sky130_fd_sc_hd__dlxbp_1 s913 (.D(net184),
    .GATE(clknet_4_3_0_clk),
    .Q(net893),
    .Q_N(net696));
 sky130_fd_sc_hd__dlxtn_2 s914 (.D(net194),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net697));
 sky130_fd_sc_hd__dlxtn_2 s915 (.D(net195),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net698));
 sky130_fd_sc_hd__dlxtn_2 s916 (.D(net203),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net904));
 sky130_fd_sc_hd__dlxtp_1 s917 (.D(net206),
    .GATE(clknet_4_3_0_clk),
    .Q(net699));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s918 (.D(net211),
    .SLEEP_B(clknet_4_2_0_clk),
    .Q(net700));
 sky130_fd_sc_hd__dfxbp_2 s919 (.CLK(clknet_4_2_0_clk),
    .D(net222),
    .Q(net702),
    .Q_N(net701));
 sky130_fd_sc_hd__dfxbp_2 s920 (.CLK(clknet_4_13_0_clk),
    .D(net248),
    .Q(net704),
    .Q_N(net703));
 sky130_fd_sc_hd__dfxtp_4 s921 (.CLK(clknet_4_13_0_clk),
    .D(net251),
    .Q(net705));
 sky130_fd_sc_hd__dfxtp_2 s922 (.CLK(clknet_4_13_0_clk),
    .D(net252),
    .Q(net706));
 sky130_fd_sc_hd__dfxtp_1 s923 (.CLK(clknet_4_13_0_clk),
    .D(net255),
    .Q(net707));
 sky130_fd_sc_hd__dlclkp_1 s924 (.CLK(clknet_4_7_0_clk),
    .GATE(net258),
    .GCLK(net708));
 sky130_fd_sc_hd__dlclkp_2 s925 (.CLK(clknet_4_12_0_clk),
    .GATE(net273),
    .GCLK(net709));
 sky130_fd_sc_hd__dlclkp_4 s926 (.CLK(clknet_4_12_0_clk),
    .GATE(net276),
    .GCLK(net875));
 sky130_fd_sc_hd__dlxbn_2 s927 (.D(net282),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net711),
    .Q_N(net710));
 sky130_fd_sc_hd__dlxbn_1 s928 (.D(net283),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net713),
    .Q_N(net712));
 sky130_fd_sc_hd__dlxbp_1 s929 (.D(net284),
    .GATE(clknet_4_6_0_clk),
    .Q(net715),
    .Q_N(net714));
 sky130_fd_sc_hd__dlxtn_2 s930 (.D(net289),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net908));
 sky130_fd_sc_hd__dlxtn_1 s931 (.D(net290),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net716));
 sky130_fd_sc_hd__dlxtn_4 s932 (.D(net294),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net717));
 sky130_fd_sc_hd__dlxtp_1 s933 (.D(net297),
    .GATE(clknet_4_6_0_clk),
    .Q(net718));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s934 (.D(net301),
    .SLEEP_B(clknet_4_6_0_clk),
    .Q(net719));
 sky130_fd_sc_hd__dfxbp_1 s935 (.CLK(clknet_4_3_0_clk),
    .D(net308),
    .Q(net721),
    .Q_N(net720));
 sky130_fd_sc_hd__dfxbp_1 s936 (.CLK(clknet_4_3_0_clk),
    .D(net313),
    .Q(net883),
    .Q_N(net722));
 sky130_fd_sc_hd__dfxtp_2 s937 (.CLK(clknet_4_8_0_clk),
    .D(net317),
    .Q(net723));
 sky130_fd_sc_hd__dfxtp_1 s938 (.CLK(clknet_4_13_0_clk),
    .D(net345),
    .Q(net724));
 sky130_fd_sc_hd__dfxtp_2 s939 (.CLK(clknet_4_13_0_clk),
    .D(net351),
    .Q(net725));
 sky130_fd_sc_hd__dlclkp_1 s940 (.CLK(clknet_4_13_0_clk),
    .GATE(net356),
    .GCLK(net726));
 sky130_fd_sc_hd__dlclkp_2 s941 (.CLK(clknet_4_13_0_clk),
    .GATE(net360),
    .GCLK(net727));
 sky130_fd_sc_hd__dlclkp_4 s942 (.CLK(clknet_4_13_0_clk),
    .GATE(net362),
    .GCLK(net728));
 sky130_fd_sc_hd__dlxbn_1 s943 (.D(net366),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net730),
    .Q_N(net729));
 sky130_fd_sc_hd__dlxbn_1 s944 (.D(net367),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net732),
    .Q_N(net731));
 sky130_fd_sc_hd__dlxbp_1 s945 (.D(net372),
    .GATE(clknet_4_12_0_clk),
    .Q(net734),
    .Q_N(net733));
 sky130_fd_sc_hd__dlxtn_2 s946 (.D(net375),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net735));
 sky130_fd_sc_hd__dlxtn_4 s947 (.D(net379),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net736));
 sky130_fd_sc_hd__dlxtn_1 s948 (.D(net380),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net737));
 sky130_fd_sc_hd__dlxtp_1 s949 (.D(net385),
    .GATE(clknet_4_12_0_clk),
    .Q(net738));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s950 (.D(net389),
    .SLEEP_B(clknet_4_9_0_clk),
    .Q(net739));
 sky130_fd_sc_hd__dfxbp_1 s951 (.CLK(clknet_4_9_0_clk),
    .D(net390),
    .Q(net741),
    .Q_N(net740));
 sky130_fd_sc_hd__dfxbp_1 s952 (.CLK(clknet_4_14_0_clk),
    .D(net397),
    .Q(net743),
    .Q_N(net742));
 sky130_fd_sc_hd__dfxtp_1 s953 (.CLK(clknet_4_8_0_clk),
    .D(net399),
    .Q(net866));
 sky130_fd_sc_hd__dfxtp_2 s954 (.CLK(clknet_4_14_0_clk),
    .D(net401),
    .Q(net744));
 sky130_fd_sc_hd__dfxtp_2 s955 (.CLK(clknet_4_8_0_clk),
    .D(net410),
    .Q(net745));
 sky130_fd_sc_hd__dlclkp_1 s956 (.CLK(clknet_4_9_0_clk),
    .GATE(net411),
    .GCLK(net746));
 sky130_fd_sc_hd__dlclkp_2 s957 (.CLK(clknet_4_8_0_clk),
    .GATE(net420),
    .GCLK(net891));
 sky130_fd_sc_hd__dlclkp_4 s958 (.CLK(clknet_4_8_0_clk),
    .GATE(net428),
    .GCLK(net879));
 sky130_fd_sc_hd__dlxbn_1 s959 (.D(net430),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net748),
    .Q_N(net747));
 sky130_fd_sc_hd__dlxbn_1 s960 (.D(net432),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net750),
    .Q_N(net749));
 sky130_fd_sc_hd__dlxbp_1 s961 (.D(net434),
    .GATE(clknet_4_8_0_clk),
    .Q(net752),
    .Q_N(net751));
 sky130_fd_sc_hd__dlxtn_2 s962 (.D(net459),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net753));
 sky130_fd_sc_hd__dlxtn_1 s963 (.D(net465),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net754));
 sky130_fd_sc_hd__dlxtn_1 s964 (.D(net467),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net755));
 sky130_fd_sc_hd__dlxtp_1 s965 (.D(net473),
    .GATE(clknet_4_15_0_clk),
    .Q(net756));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s966 (.D(net475),
    .SLEEP_B(clknet_4_14_0_clk),
    .Q(net757));
 sky130_fd_sc_hd__dfxbp_1 s967 (.CLK(clknet_4_14_0_clk),
    .D(net479),
    .Q(net759),
    .Q_N(net758));
 sky130_fd_sc_hd__dfxbp_2 s968 (.CLK(clknet_4_15_0_clk),
    .D(net483),
    .Q(net761),
    .Q_N(net760));
 sky130_fd_sc_hd__dfxtp_2 s969 (.CLK(clknet_4_14_0_clk),
    .D(net494),
    .Q(net762));
 sky130_fd_sc_hd__dfxtp_2 s970 (.CLK(clknet_4_11_0_clk),
    .D(net503),
    .Q(net763));
 sky130_fd_sc_hd__dfxtp_1 s971 (.CLK(clknet_4_14_0_clk),
    .D(net505),
    .Q(net874));
 sky130_fd_sc_hd__dlclkp_1 s972 (.CLK(clknet_4_11_0_clk),
    .GATE(net514),
    .GCLK(net764));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(in0),
    .X(net765));
 sky130_fd_sc_hd__buf_1 input2 (.A(in1),
    .X(net766));
 sky130_fd_sc_hd__buf_2 input3 (.A(in10),
    .X(net767));
 sky130_fd_sc_hd__buf_2 input4 (.A(in11),
    .X(net768));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(in12),
    .X(net769));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(in13),
    .X(net770));
 sky130_fd_sc_hd__buf_4 input7 (.A(in14),
    .X(net771));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(in15),
    .X(net772));
 sky130_fd_sc_hd__buf_1 input9 (.A(in16),
    .X(net773));
 sky130_fd_sc_hd__buf_2 input10 (.A(in17),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(in18),
    .X(net775));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(in19),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(in2),
    .X(net777));
 sky130_fd_sc_hd__buf_2 input14 (.A(in20),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(in21),
    .X(net779));
 sky130_fd_sc_hd__buf_2 input16 (.A(in22),
    .X(net780));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(in23),
    .X(net781));
 sky130_fd_sc_hd__buf_1 input18 (.A(in24),
    .X(net782));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(in25),
    .X(net783));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(in26),
    .X(net784));
 sky130_fd_sc_hd__buf_2 input21 (.A(in27),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(in28),
    .X(net786));
 sky130_fd_sc_hd__clkbuf_4 input23 (.A(in29),
    .X(net787));
 sky130_fd_sc_hd__buf_12 input24 (.A(in3),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(in30),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_4 input26 (.A(in31),
    .X(net790));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(in32),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(in33),
    .X(net792));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(in34),
    .X(net793));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(in35),
    .X(net794));
 sky130_fd_sc_hd__buf_2 input31 (.A(in36),
    .X(net795));
 sky130_fd_sc_hd__buf_1 input32 (.A(in37),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(in38),
    .X(net797));
 sky130_fd_sc_hd__buf_2 input34 (.A(in39),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_4 input35 (.A(in4),
    .X(net799));
 sky130_fd_sc_hd__buf_6 input36 (.A(in40),
    .X(net800));
 sky130_fd_sc_hd__buf_4 input37 (.A(in41),
    .X(net801));
 sky130_fd_sc_hd__buf_2 input38 (.A(in42),
    .X(net802));
 sky130_fd_sc_hd__buf_4 input39 (.A(in43),
    .X(net803));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(in44),
    .X(net804));
 sky130_fd_sc_hd__buf_4 input41 (.A(in45),
    .X(net805));
 sky130_fd_sc_hd__buf_2 input42 (.A(in46),
    .X(net806));
 sky130_fd_sc_hd__buf_1 input43 (.A(in47),
    .X(net807));
 sky130_fd_sc_hd__clkbuf_4 input44 (.A(in48),
    .X(net808));
 sky130_fd_sc_hd__buf_1 input45 (.A(in49),
    .X(net809));
 sky130_fd_sc_hd__buf_1 input46 (.A(in5),
    .X(net810));
 sky130_fd_sc_hd__dlymetal6s2s_1 input47 (.A(in50),
    .X(net811));
 sky130_fd_sc_hd__buf_2 input48 (.A(in51),
    .X(net812));
 sky130_fd_sc_hd__buf_2 input49 (.A(in52),
    .X(net813));
 sky130_fd_sc_hd__buf_2 input50 (.A(in53),
    .X(net814));
 sky130_fd_sc_hd__dlymetal6s2s_1 input51 (.A(in54),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(in55),
    .X(net816));
 sky130_fd_sc_hd__buf_4 input53 (.A(in56),
    .X(net817));
 sky130_fd_sc_hd__buf_2 input54 (.A(in57),
    .X(net818));
 sky130_fd_sc_hd__buf_4 input55 (.A(in58),
    .X(net819));
 sky130_fd_sc_hd__buf_1 input56 (.A(in59),
    .X(net820));
 sky130_fd_sc_hd__dlymetal6s2s_1 input57 (.A(in6),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(in60),
    .X(net822));
 sky130_fd_sc_hd__buf_2 input59 (.A(in61),
    .X(net823));
 sky130_fd_sc_hd__buf_4 input60 (.A(in62),
    .X(net824));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(in63),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(in64),
    .X(net826));
 sky130_fd_sc_hd__buf_1 input63 (.A(in65),
    .X(net827));
 sky130_fd_sc_hd__buf_1 input64 (.A(in66),
    .X(net828));
 sky130_fd_sc_hd__buf_1 input65 (.A(in67),
    .X(net829));
 sky130_fd_sc_hd__buf_1 input66 (.A(in68),
    .X(net830));
 sky130_fd_sc_hd__clkbuf_4 input67 (.A(in69),
    .X(net831));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(in7),
    .X(net832));
 sky130_fd_sc_hd__clkbuf_4 input69 (.A(in70),
    .X(net833));
 sky130_fd_sc_hd__buf_1 input70 (.A(in71),
    .X(net834));
 sky130_fd_sc_hd__buf_2 input71 (.A(in72),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_2 input72 (.A(in73),
    .X(net836));
 sky130_fd_sc_hd__clkbuf_4 input73 (.A(in74),
    .X(net837));
 sky130_fd_sc_hd__buf_2 input74 (.A(in75),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_2 input75 (.A(in76),
    .X(net839));
 sky130_fd_sc_hd__buf_1 input76 (.A(in77),
    .X(net840));
 sky130_fd_sc_hd__buf_1 input77 (.A(in78),
    .X(net841));
 sky130_fd_sc_hd__buf_1 input78 (.A(in79),
    .X(net842));
 sky130_fd_sc_hd__buf_1 input79 (.A(in8),
    .X(net843));
 sky130_fd_sc_hd__buf_1 input80 (.A(in80),
    .X(net844));
 sky130_fd_sc_hd__buf_1 input81 (.A(in81),
    .X(net845));
 sky130_fd_sc_hd__clkbuf_4 input82 (.A(in82),
    .X(net846));
 sky130_fd_sc_hd__buf_2 input83 (.A(in83),
    .X(net847));
 sky130_fd_sc_hd__buf_1 input84 (.A(in84),
    .X(net848));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(in85),
    .X(net849));
 sky130_fd_sc_hd__buf_1 input86 (.A(in86),
    .X(net850));
 sky130_fd_sc_hd__buf_1 input87 (.A(in87),
    .X(net851));
 sky130_fd_sc_hd__buf_1 input88 (.A(in88),
    .X(net852));
 sky130_fd_sc_hd__buf_1 input89 (.A(in89),
    .X(net853));
 sky130_fd_sc_hd__buf_4 input90 (.A(in9),
    .X(net854));
 sky130_fd_sc_hd__buf_1 input91 (.A(in90),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_4 input92 (.A(in91),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_4 input93 (.A(in92),
    .X(net857));
 sky130_fd_sc_hd__buf_4 input94 (.A(in93),
    .X(net858));
 sky130_fd_sc_hd__buf_2 input95 (.A(in94),
    .X(net859));
 sky130_fd_sc_hd__buf_1 input96 (.A(in95),
    .X(net860));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(in96),
    .X(net861));
 sky130_fd_sc_hd__buf_2 input98 (.A(in97),
    .X(net862));
 sky130_fd_sc_hd__clkbuf_2 input99 (.A(in98),
    .X(net863));
 sky130_fd_sc_hd__buf_1 input100 (.A(in99),
    .X(net864));
 sky130_fd_sc_hd__buf_2 output101 (.A(net983),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output102 (.A(net866),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output103 (.A(net867),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_1 output104 (.A(clknet_1_1__leaf_net868),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output105 (.A(net985),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output106 (.A(net870),
    .X(out14));
 sky130_fd_sc_hd__clkbuf_4 output107 (.A(net871),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output108 (.A(net1088),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output109 (.A(net873),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output110 (.A(net874),
    .X(out2));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(clknet_1_0__leaf_net875),
    .X(out20));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(net876),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output113 (.A(net877),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(clknet_1_1__leaf_net878),
    .X(out23));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(clknet_1_0__leaf_net879),
    .X(out24));
 sky130_fd_sc_hd__clkbuf_1 output116 (.A(clknet_1_1__leaf_net880),
    .X(out25));
 sky130_fd_sc_hd__buf_2 output117 (.A(net968),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output118 (.A(net882),
    .X(out27));
 sky130_fd_sc_hd__buf_2 output119 (.A(net883),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output120 (.A(net884),
    .X(out29));
 sky130_fd_sc_hd__buf_2 output121 (.A(net885),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output122 (.A(net886),
    .X(out31));
 sky130_fd_sc_hd__clkbuf_1 output123 (.A(clknet_1_1__leaf_net887),
    .X(out32));
 sky130_fd_sc_hd__buf_2 output124 (.A(net888),
    .X(out33));
 sky130_fd_sc_hd__clkbuf_4 output125 (.A(net889),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output126 (.A(net890),
    .X(out35));
 sky130_fd_sc_hd__clkbuf_1 output127 (.A(clknet_1_1__leaf_net891),
    .X(out37));
 sky130_fd_sc_hd__clkbuf_1 output128 (.A(clknet_1_1__leaf_net892),
    .X(out38));
 sky130_fd_sc_hd__buf_2 output129 (.A(net893),
    .X(out39));
 sky130_fd_sc_hd__clkbuf_1 output130 (.A(clknet_1_0__leaf_net894),
    .X(out43));
 sky130_fd_sc_hd__clkbuf_1 output131 (.A(net895),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output132 (.A(net896),
    .X(out46));
 sky130_fd_sc_hd__buf_2 output133 (.A(net897),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output134 (.A(net898),
    .X(out48));
 sky130_fd_sc_hd__buf_2 output135 (.A(net899),
    .X(out49));
 sky130_fd_sc_hd__buf_2 output136 (.A(net900),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output137 (.A(net901),
    .X(out51));
 sky130_fd_sc_hd__buf_2 output138 (.A(net902),
    .X(out52));
 sky130_fd_sc_hd__clkbuf_4 output139 (.A(net903),
    .X(out53));
 sky130_fd_sc_hd__buf_2 output140 (.A(net904),
    .X(out54));
 sky130_fd_sc_hd__buf_2 output141 (.A(net905),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output142 (.A(net906),
    .X(out57));
 sky130_fd_sc_hd__clkbuf_1 output143 (.A(clknet_1_0__leaf_net907),
    .X(out58));
 sky130_fd_sc_hd__buf_2 output144 (.A(net908),
    .X(out59));
 sky130_fd_sc_hd__clkbuf_1 output145 (.A(clknet_1_1__leaf_net909),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_1 output146 (.A(clknet_1_0__leaf_net910),
    .X(out60));
 sky130_fd_sc_hd__clkbuf_1 output147 (.A(clknet_1_0__leaf_net911),
    .X(out62));
 sky130_fd_sc_hd__clkbuf_1 output148 (.A(clknet_1_0__leaf_net912),
    .X(out63));
 sky130_fd_sc_hd__buf_2 output149 (.A(net913),
    .X(out64));
 sky130_fd_sc_hd__buf_2 output150 (.A(net914),
    .X(out66));
 sky130_fd_sc_hd__buf_2 output151 (.A(net915),
    .X(out67));
 sky130_fd_sc_hd__buf_2 output152 (.A(net916),
    .X(out68));
 sky130_fd_sc_hd__clkbuf_1 output153 (.A(net917),
    .X(out69));
 sky130_fd_sc_hd__buf_2 output154 (.A(net918),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output155 (.A(net919),
    .X(out70));
 sky130_fd_sc_hd__buf_2 output156 (.A(net920),
    .X(out71));
 sky130_fd_sc_hd__buf_2 output157 (.A(net921),
    .X(out74));
 sky130_fd_sc_hd__clkbuf_1 output158 (.A(clknet_1_0__leaf_net922),
    .X(out75));
 sky130_fd_sc_hd__buf_2 output159 (.A(net923),
    .X(out76));
 sky130_fd_sc_hd__buf_2 output160 (.A(net924),
    .X(out78));
 sky130_fd_sc_hd__clkbuf_1 output161 (.A(clknet_1_0__leaf_net925),
    .X(out79));
 sky130_fd_sc_hd__buf_2 output162 (.A(net926),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output163 (.A(net927),
    .X(out80));
 sky130_fd_sc_hd__clkbuf_4 output164 (.A(net928),
    .X(out81));
 sky130_fd_sc_hd__buf_2 output165 (.A(net929),
    .X(out82));
 sky130_fd_sc_hd__buf_2 output166 (.A(net930),
    .X(out84));
 sky130_fd_sc_hd__buf_2 output167 (.A(net931),
    .X(out85));
 sky130_fd_sc_hd__buf_2 output168 (.A(net932),
    .X(out86));
 sky130_fd_sc_hd__buf_2 output169 (.A(net933),
    .X(out87));
 sky130_fd_sc_hd__buf_2 output170 (.A(net934),
    .X(out88));
 sky130_fd_sc_hd__buf_2 output171 (.A(net998),
    .X(out89));
 sky130_fd_sc_hd__buf_2 output172 (.A(net936),
    .X(out9));
 sky130_fd_sc_hd__buf_2 output173 (.A(net937),
    .X(out90));
 sky130_fd_sc_hd__buf_2 output174 (.A(net938),
    .X(out91));
 sky130_fd_sc_hd__buf_2 output175 (.A(net939),
    .X(out93));
 sky130_fd_sc_hd__buf_2 output176 (.A(net940),
    .X(out94));
 sky130_fd_sc_hd__buf_2 output177 (.A(net941),
    .X(out95));
 sky130_fd_sc_hd__buf_2 output178 (.A(net942),
    .X(out96));
 sky130_fd_sc_hd__buf_2 output179 (.A(net943),
    .X(out97));
 sky130_fd_sc_hd__clkbuf_1 output180 (.A(net944),
    .X(out98));
 sky130_fd_sc_hd__buf_2 output181 (.A(net945),
    .X(out99));
 sky130_fd_sc_hd__buf_4 fanout182 (.A(net43),
    .X(net946));
 sky130_fd_sc_hd__clkbuf_4 fanout183 (.A(net253),
    .X(net947));
 sky130_fd_sc_hd__buf_4 fanout184 (.A(net242),
    .X(net948));
 sky130_fd_sc_hd__buf_2 fanout185 (.A(net950),
    .X(net949));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout186 (.A(net951),
    .X(net950));
 sky130_fd_sc_hd__clkbuf_4 fanout187 (.A(net952),
    .X(net951));
 sky130_fd_sc_hd__clkbuf_4 fanout188 (.A(net123),
    .X(net952));
 sky130_fd_sc_hd__clkbuf_4 fanout189 (.A(net85),
    .X(net953));
 sky130_fd_sc_hd__clkbuf_4 fanout190 (.A(net41),
    .X(net954));
 sky130_fd_sc_hd__buf_2 fanout191 (.A(net956),
    .X(net955));
 sky130_fd_sc_hd__clkbuf_2 fanout192 (.A(net957),
    .X(net956));
 sky130_fd_sc_hd__buf_2 fanout193 (.A(net958),
    .X(net957));
 sky130_fd_sc_hd__clkbuf_4 fanout194 (.A(net118),
    .X(net958));
 sky130_fd_sc_hd__clkbuf_4 fanout195 (.A(net40),
    .X(net959));
 sky130_fd_sc_hd__buf_4 fanout196 (.A(net39),
    .X(net960));
 sky130_fd_sc_hd__buf_4 fanout197 (.A(net32),
    .X(net961));
 sky130_fd_sc_hd__buf_2 fanout198 (.A(net32),
    .X(net962));
 sky130_fd_sc_hd__buf_4 fanout199 (.A(net913),
    .X(net963));
 sky130_fd_sc_hd__buf_12 fanout200 (.A(net31),
    .X(net964));
 sky130_fd_sc_hd__clkbuf_2 fanout201 (.A(net1039),
    .X(net965));
 sky130_fd_sc_hd__buf_4 fanout202 (.A(net967),
    .X(net966));
 sky130_fd_sc_hd__clkbuf_4 fanout203 (.A(net37),
    .X(net967));
 sky130_fd_sc_hd__buf_8 fanout204 (.A(net881),
    .X(net968));
 sky130_fd_sc_hd__buf_12 fanout205 (.A(net30),
    .X(net969));
 sky130_fd_sc_hd__buf_4 fanout206 (.A(net35),
    .X(net970));
 sky130_fd_sc_hd__buf_8 fanout207 (.A(net29),
    .X(net971));
 sky130_fd_sc_hd__buf_8 fanout208 (.A(net27),
    .X(net972));
 sky130_fd_sc_hd__buf_6 fanout209 (.A(net974),
    .X(net973));
 sky130_fd_sc_hd__buf_8 fanout210 (.A(net871),
    .X(net974));
 sky130_fd_sc_hd__buf_12 fanout211 (.A(net28),
    .X(net975));
 sky130_fd_sc_hd__buf_12 fanout212 (.A(net23),
    .X(net976));
 sky130_fd_sc_hd__clkbuf_4 fanout213 (.A(net978),
    .X(net977));
 sky130_fd_sc_hd__buf_12 fanout214 (.A(net979),
    .X(net978));
 sky130_fd_sc_hd__buf_8 fanout215 (.A(net21),
    .X(net979));
 sky130_fd_sc_hd__buf_12 fanout216 (.A(net20),
    .X(net980));
 sky130_fd_sc_hd__buf_2 fanout217 (.A(net20),
    .X(net981));
 sky130_fd_sc_hd__buf_12 fanout218 (.A(net865),
    .X(net982));
 sky130_fd_sc_hd__buf_2 fanout219 (.A(net1058),
    .X(net983));
 sky130_fd_sc_hd__buf_2 fanout220 (.A(net985),
    .X(net984));
 sky130_fd_sc_hd__clkbuf_4 fanout221 (.A(net869),
    .X(net985));
 sky130_fd_sc_hd__buf_12 fanout222 (.A(net19),
    .X(net986));
 sky130_fd_sc_hd__buf_8 fanout223 (.A(net16),
    .X(net987));
 sky130_fd_sc_hd__buf_2 max_cap224 (.A(net719),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_4 wire225 (.A(net699),
    .X(net989));
 sky130_fd_sc_hd__buf_4 max_cap226 (.A(net682),
    .X(net990));
 sky130_fd_sc_hd__clkbuf_8 fanout227 (.A(net681),
    .X(net991));
 sky130_fd_sc_hd__buf_4 fanout228 (.A(net680),
    .X(net992));
 sky130_fd_sc_hd__clkbuf_4 fanout229 (.A(net994),
    .X(net993));
 sky130_fd_sc_hd__clkbuf_2 fanout230 (.A(net995),
    .X(net994));
 sky130_fd_sc_hd__clkbuf_4 fanout231 (.A(net668),
    .X(net995));
 sky130_fd_sc_hd__buf_4 fanout232 (.A(net133),
    .X(net996));
 sky130_fd_sc_hd__clkbuf_4 fanout233 (.A(net134),
    .X(net997));
 sky130_fd_sc_hd__buf_12 fanout234 (.A(net935),
    .X(net998));
 sky130_fd_sc_hd__buf_12 fanout235 (.A(net854),
    .X(net999));
 sky130_fd_sc_hd__clkbuf_4 fanout236 (.A(net773),
    .X(net1000));
 sky130_fd_sc_hd__buf_12 fanout237 (.A(net772),
    .X(net1001));
 sky130_fd_sc_hd__clkbuf_2 fanout238 (.A(net772),
    .X(net1002));
 sky130_fd_sc_hd__buf_4 fanout239 (.A(net1004),
    .X(net1003));
 sky130_fd_sc_hd__buf_4 fanout240 (.A(net843),
    .X(net1004));
 sky130_fd_sc_hd__buf_12 fanout241 (.A(net771),
    .X(net1005));
 sky130_fd_sc_hd__buf_4 fanout242 (.A(net1007),
    .X(net1006));
 sky130_fd_sc_hd__clkbuf_4 fanout243 (.A(net832),
    .X(net1007));
 sky130_fd_sc_hd__buf_4 fanout244 (.A(net821),
    .X(net1008));
 sky130_fd_sc_hd__buf_2 fanout245 (.A(net821),
    .X(net1009));
 sky130_fd_sc_hd__buf_4 fanout246 (.A(net769),
    .X(net1010));
 sky130_fd_sc_hd__buf_2 fanout247 (.A(net769),
    .X(net1011));
 sky130_fd_sc_hd__buf_4 fanout248 (.A(net810),
    .X(net1012));
 sky130_fd_sc_hd__buf_4 fanout249 (.A(net768),
    .X(net1013));
 sky130_fd_sc_hd__buf_12 fanout250 (.A(net799),
    .X(net1014));
 sky130_fd_sc_hd__buf_4 fanout251 (.A(net796),
    .X(net1015));
 sky130_fd_sc_hd__clkbuf_8 fanout252 (.A(net789),
    .X(net1016));
 sky130_fd_sc_hd__clkbuf_4 fanout253 (.A(net1018),
    .X(net1017));
 sky130_fd_sc_hd__clkbuf_4 fanout254 (.A(net788),
    .X(net1018));
 sky130_fd_sc_hd__buf_12 fanout255 (.A(net1020),
    .X(net1019));
 sky130_fd_sc_hd__buf_12 fanout256 (.A(net788),
    .X(net1020));
 sky130_fd_sc_hd__buf_4 fanout257 (.A(net1022),
    .X(net1021));
 sky130_fd_sc_hd__clkbuf_4 fanout258 (.A(net788),
    .X(net1022));
 sky130_fd_sc_hd__buf_4 fanout259 (.A(net766),
    .X(net1023));
 sky130_fd_sc_hd__buf_4 fanout260 (.A(net783),
    .X(net1024));
 sky130_fd_sc_hd__clkbuf_2 fanout261 (.A(net783),
    .X(net1025));
 sky130_fd_sc_hd__buf_4 fanout262 (.A(net782),
    .X(net1026));
 sky130_fd_sc_hd__buf_4 fanout263 (.A(net779),
    .X(net1027));
 sky130_fd_sc_hd__buf_4 fanout264 (.A(net778),
    .X(net1028));
 sky130_fd_sc_hd__clkbuf_4 fanout265 (.A(net777),
    .X(net1029));
 sky130_fd_sc_hd__buf_8 fanout266 (.A(net776),
    .X(net1030));
 sky130_fd_sc_hd__buf_12 fanout267 (.A(net775),
    .X(net1031));
 sky130_fd_sc_hd__clkbuf_8 fanout268 (.A(net774),
    .X(net1032));
 sky130_fd_sc_hd__clkbuf_8 fanout269 (.A(net765),
    .X(net1033));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net764 (.A(net764),
    .X(clknet_0_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net764 (.A(clknet_0_net764),
    .X(clknet_1_0__leaf_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net764 (.A(clknet_0_net764),
    .X(clknet_1_1__leaf_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net650 (.A(net650),
    .X(clknet_0_net650));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net650 (.A(clknet_0_net650),
    .X(clknet_1_0__leaf_net650));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net650 (.A(clknet_0_net650),
    .X(clknet_1_1__leaf_net650));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net526 (.A(net526),
    .X(clknet_0_net526));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net526 (.A(clknet_0_net526),
    .X(clknet_1_0__leaf_net526));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net526 (.A(clknet_0_net526),
    .X(clknet_1_1__leaf_net526));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net527 (.A(net527),
    .X(clknet_0_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net527 (.A(clknet_0_net527),
    .X(clknet_1_0__leaf_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net527 (.A(clknet_0_net527),
    .X(clknet_1_1__leaf_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net525 (.A(net525),
    .X(clknet_0_net525));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net525 (.A(clknet_0_net525),
    .X(clknet_1_0__leaf_net525));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net525 (.A(clknet_0_net525),
    .X(clknet_1_1__leaf_net525));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net547 (.A(net547),
    .X(clknet_0_net547));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net547 (.A(clknet_0_net547),
    .X(clknet_1_0__leaf_net547));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net547 (.A(clknet_0_net547),
    .X(clknet_1_1__leaf_net547));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net879 (.A(net879),
    .X(clknet_0_net879));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net879 (.A(clknet_0_net879),
    .X(clknet_1_0__leaf_net879));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net879 (.A(clknet_0_net879),
    .X(clknet_1_1__leaf_net879));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net436 (.A(net436),
    .X(clknet_0_net436));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net436 (.A(clknet_0_net436),
    .X(clknet_1_0__leaf_net436));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net436 (.A(clknet_0_net436),
    .X(clknet_1_1__leaf_net436));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net891 (.A(net891),
    .X(clknet_0_net891));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net891 (.A(clknet_0_net891),
    .X(clknet_1_0__leaf_net891));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net891 (.A(clknet_0_net891),
    .X(clknet_1_1__leaf_net891));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net423 (.A(net423),
    .X(clknet_0_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net423 (.A(clknet_0_net423),
    .X(clknet_1_0__leaf_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net423 (.A(clknet_0_net423),
    .X(clknet_1_1__leaf_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net427 (.A(net427),
    .X(clknet_0_net427));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net427 (.A(clknet_0_net427),
    .X(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net427 (.A(clknet_0_net427),
    .X(clknet_1_1__leaf_net427));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net878 (.A(net878),
    .X(clknet_0_net878));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net878 (.A(clknet_0_net878),
    .X(clknet_1_0__leaf_net878));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net878 (.A(clknet_0_net878),
    .X(clknet_1_1__leaf_net878));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net422 (.A(net422),
    .X(clknet_0_net422));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net422 (.A(clknet_0_net422),
    .X(clknet_1_0__leaf_net422));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net422 (.A(clknet_0_net422),
    .X(clknet_1_1__leaf_net422));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net424 (.A(net424),
    .X(clknet_0_net424));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net424 (.A(clknet_0_net424),
    .X(clknet_1_0__leaf_net424));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net424 (.A(clknet_0_net424),
    .X(clknet_1_1__leaf_net424));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net746 (.A(net746),
    .X(clknet_0_net746));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net746 (.A(clknet_0_net746),
    .X(clknet_1_0__leaf_net746));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net746 (.A(clknet_0_net746),
    .X(clknet_1_1__leaf_net746));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net416 (.A(net416),
    .X(clknet_0_net416));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net416 (.A(clknet_0_net416),
    .X(clknet_1_0__leaf_net416));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net416 (.A(clknet_0_net416),
    .X(clknet_1_1__leaf_net416));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net728 (.A(net728),
    .X(clknet_0_net728));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net728 (.A(clknet_0_net728),
    .X(clknet_1_0__leaf_net728));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net728 (.A(clknet_0_net728),
    .X(clknet_1_1__leaf_net728));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net887 (.A(net887),
    .X(clknet_0_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net887 (.A(clknet_0_net887),
    .X(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net887 (.A(clknet_0_net887),
    .X(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net365 (.A(net365),
    .X(clknet_0_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net365 (.A(clknet_0_net365),
    .X(clknet_1_0__leaf_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net365 (.A(clknet_0_net365),
    .X(clknet_1_1__leaf_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net496 (.A(net496),
    .X(clknet_0_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net496 (.A(clknet_0_net496),
    .X(clknet_1_0__leaf_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net496 (.A(clknet_0_net496),
    .X(clknet_1_1__leaf_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net727 (.A(net727),
    .X(clknet_0_net727));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net727 (.A(clknet_0_net727),
    .X(clknet_1_0__leaf_net727));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net727 (.A(clknet_0_net727),
    .X(clknet_1_1__leaf_net727));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net466 (.A(net466),
    .X(clknet_0_net466));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net466 (.A(clknet_0_net466),
    .X(clknet_1_0__leaf_net466));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net466 (.A(clknet_0_net466),
    .X(clknet_1_1__leaf_net466));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net484 (.A(net484),
    .X(clknet_0_net484));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net484 (.A(clknet_0_net484),
    .X(clknet_1_0__leaf_net484));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net484 (.A(clknet_0_net484),
    .X(clknet_1_1__leaf_net484));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net368 (.A(net368),
    .X(clknet_0_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net368 (.A(clknet_0_net368),
    .X(clknet_1_0__leaf_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net368 (.A(clknet_0_net368),
    .X(clknet_1_1__leaf_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net376 (.A(net376),
    .X(clknet_0_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net376 (.A(clknet_0_net376),
    .X(clknet_1_0__leaf_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net376 (.A(clknet_0_net376),
    .X(clknet_1_1__leaf_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net364 (.A(net364),
    .X(clknet_0_net364));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net364 (.A(clknet_0_net364),
    .X(clknet_1_0__leaf_net364));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net364 (.A(clknet_0_net364),
    .X(clknet_1_1__leaf_net364));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net382 (.A(net382),
    .X(clknet_0_net382));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net382 (.A(clknet_0_net382),
    .X(clknet_1_0__leaf_net382));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net382 (.A(clknet_0_net382),
    .X(clknet_1_1__leaf_net382));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net398 (.A(net398),
    .X(clknet_0_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_0__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_1__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net384 (.A(net384),
    .X(clknet_0_net384));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net384 (.A(clknet_0_net384),
    .X(clknet_1_0__leaf_net384));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net384 (.A(clknet_0_net384),
    .X(clknet_1_1__leaf_net384));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net363 (.A(net363),
    .X(clknet_0_net363));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net363 (.A(clknet_0_net363),
    .X(clknet_1_0__leaf_net363));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net363 (.A(clknet_0_net363),
    .X(clknet_1_1__leaf_net363));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net361 (.A(net361),
    .X(clknet_0_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net361 (.A(clknet_0_net361),
    .X(clknet_1_0__leaf_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net361 (.A(clknet_0_net361),
    .X(clknet_1_1__leaf_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net726 (.A(net726),
    .X(clknet_0_net726));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net726 (.A(clknet_0_net726),
    .X(clknet_1_0__leaf_net726));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net726 (.A(clknet_0_net726),
    .X(clknet_1_1__leaf_net726));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net396 (.A(net396),
    .X(clknet_0_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_0__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_1__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net506 (.A(net506),
    .X(clknet_0_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net506 (.A(clknet_0_net506),
    .X(clknet_1_0__leaf_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net506 (.A(clknet_0_net506),
    .X(clknet_1_1__leaf_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net532 (.A(net532),
    .X(clknet_0_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net532 (.A(clknet_0_net532),
    .X(clknet_1_0__leaf_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net532 (.A(clknet_0_net532),
    .X(clknet_1_1__leaf_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net499 (.A(net499),
    .X(clknet_0_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net499 (.A(clknet_0_net499),
    .X(clknet_1_0__leaf_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net499 (.A(clknet_0_net499),
    .X(clknet_1_1__leaf_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net875 (.A(net875),
    .X(clknet_0_net875));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net875 (.A(clknet_0_net875),
    .X(clknet_1_0__leaf_net875));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net875 (.A(clknet_0_net875),
    .X(clknet_1_1__leaf_net875));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net383 (.A(net383),
    .X(clknet_0_net383));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net383 (.A(clknet_0_net383),
    .X(clknet_1_0__leaf_net383));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net383 (.A(clknet_0_net383),
    .X(clknet_1_1__leaf_net383));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net278 (.A(net278),
    .X(clknet_0_net278));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net278 (.A(clknet_0_net278),
    .X(clknet_1_0__leaf_net278));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net278 (.A(clknet_0_net278),
    .X(clknet_1_1__leaf_net278));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net300 (.A(net300),
    .X(clknet_0_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net300 (.A(clknet_0_net300),
    .X(clknet_1_0__leaf_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net300 (.A(clknet_0_net300),
    .X(clknet_1_1__leaf_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net293 (.A(net293),
    .X(clknet_0_net293));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net293 (.A(clknet_0_net293),
    .X(clknet_1_0__leaf_net293));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net293 (.A(clknet_0_net293),
    .X(clknet_1_1__leaf_net293));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net314 (.A(net314),
    .X(clknet_0_net314));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net314 (.A(net1059),
    .X(clknet_1_0__leaf_net314));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net314 (.A(clknet_0_net314),
    .X(clknet_1_1__leaf_net314));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net316 (.A(net316),
    .X(clknet_0_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net316 (.A(clknet_0_net316),
    .X(clknet_1_0__leaf_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net316 (.A(clknet_0_net316),
    .X(clknet_1_1__leaf_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net303 (.A(net303),
    .X(clknet_0_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net303 (.A(clknet_0_net303),
    .X(clknet_1_0__leaf_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net303 (.A(clknet_0_net303),
    .X(clknet_1_1__leaf_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net912 (.A(net912),
    .X(clknet_0_net912));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net912 (.A(clknet_0_net912),
    .X(clknet_1_0__leaf_net912));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net912 (.A(clknet_0_net912),
    .X(clknet_1_1__leaf_net912));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net277 (.A(net277),
    .X(clknet_0_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net277 (.A(clknet_0_net277),
    .X(clknet_1_0__leaf_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net277 (.A(clknet_0_net277),
    .X(clknet_1_1__leaf_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net709 (.A(net709),
    .X(clknet_0_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net709 (.A(clknet_0_net709),
    .X(clknet_1_0__leaf_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net709 (.A(clknet_0_net709),
    .X(clknet_1_1__leaf_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net489 (.A(net489),
    .X(clknet_0_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_0__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_1__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net478 (.A(net478),
    .X(clknet_0_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net478 (.A(clknet_0_net478),
    .X(clknet_1_0__leaf_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net478 (.A(clknet_0_net478),
    .X(clknet_1_1__leaf_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net275 (.A(net275),
    .X(clknet_0_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net275 (.A(clknet_0_net275),
    .X(clknet_1_0__leaf_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net275 (.A(clknet_0_net275),
    .X(clknet_1_1__leaf_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net708 (.A(net708),
    .X(clknet_0_net708));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net708 (.A(clknet_0_net708),
    .X(clknet_1_0__leaf_net708));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net708 (.A(clknet_0_net708),
    .X(clknet_1_1__leaf_net708));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net335 (.A(net335),
    .X(clknet_0_net335));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net335 (.A(clknet_0_net335),
    .X(clknet_1_0__leaf_net335));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net335 (.A(clknet_0_net335),
    .X(clknet_1_1__leaf_net335));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net907 (.A(net907),
    .X(clknet_0_net907));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net907 (.A(clknet_0_net907),
    .X(clknet_1_0__leaf_net907));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net907 (.A(clknet_0_net907),
    .X(clknet_1_1__leaf_net907));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net894 (.A(net894),
    .X(clknet_0_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net894 (.A(clknet_0_net894),
    .X(clknet_1_0__leaf_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net894 (.A(clknet_0_net894),
    .X(clknet_1_1__leaf_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net330 (.A(net330),
    .X(clknet_0_net330));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net330 (.A(clknet_0_net330),
    .X(clknet_1_0__leaf_net330));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net330 (.A(clknet_0_net330),
    .X(clknet_1_1__leaf_net330));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net339 (.A(net339),
    .X(clknet_0_net339));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net339 (.A(clknet_0_net339),
    .X(clknet_1_0__leaf_net339));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net339 (.A(clknet_0_net339),
    .X(clknet_1_1__leaf_net339));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net338 (.A(net338),
    .X(clknet_0_net338));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net338 (.A(clknet_0_net338),
    .X(clknet_1_0__leaf_net338));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net338 (.A(clknet_0_net338),
    .X(clknet_1_1__leaf_net338));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net262 (.A(net262),
    .X(clknet_0_net262));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net262 (.A(clknet_0_net262),
    .X(clknet_1_0__leaf_net262));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net262 (.A(clknet_0_net262),
    .X(clknet_1_1__leaf_net262));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net265 (.A(net265),
    .X(clknet_0_net265));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net265 (.A(clknet_0_net265),
    .X(clknet_1_0__leaf_net265));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net265 (.A(clknet_0_net265),
    .X(clknet_1_1__leaf_net265));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net259 (.A(net259),
    .X(clknet_0_net259));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net259 (.A(clknet_0_net259),
    .X(clknet_1_0__leaf_net259));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net259 (.A(clknet_0_net259),
    .X(clknet_1_1__leaf_net259));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net691 (.A(net691),
    .X(clknet_0_net691));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net691 (.A(clknet_0_net691),
    .X(clknet_1_0__leaf_net691));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net691 (.A(clknet_0_net691),
    .X(clknet_1_1__leaf_net691));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net185 (.A(net185),
    .X(clknet_0_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net185 (.A(clknet_0_net185),
    .X(clknet_1_0__leaf_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net185 (.A(clknet_0_net185),
    .X(clknet_1_1__leaf_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net868 (.A(net868),
    .X(clknet_0_net868));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net868 (.A(clknet_0_net868),
    .X(clknet_1_0__leaf_net868));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net868 (.A(clknet_0_net868),
    .X(clknet_1_1__leaf_net868));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net311 (.A(net311),
    .X(clknet_0_net311));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net311 (.A(clknet_0_net311),
    .X(clknet_1_0__leaf_net311));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net311 (.A(clknet_0_net311),
    .X(clknet_1_1__leaf_net311));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net287 (.A(net287),
    .X(clknet_0_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net287 (.A(clknet_0_net287),
    .X(clknet_1_0__leaf_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net287 (.A(clknet_0_net287),
    .X(clknet_1_1__leaf_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net911 (.A(net911),
    .X(clknet_0_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net911 (.A(clknet_0_net911),
    .X(clknet_1_0__leaf_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net911 (.A(clknet_0_net911),
    .X(clknet_1_1__leaf_net911));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net306 (.A(net306),
    .X(clknet_0_net306));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net306 (.A(clknet_0_net306),
    .X(clknet_1_0__leaf_net306));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net306 (.A(clknet_0_net306),
    .X(clknet_1_1__leaf_net306));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net909 (.A(net909),
    .X(clknet_0_net909));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net909 (.A(clknet_0_net909),
    .X(clknet_1_0__leaf_net909));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net909 (.A(clknet_0_net909),
    .X(clknet_1_1__leaf_net909));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net307 (.A(net307),
    .X(clknet_0_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net307 (.A(clknet_0_net307),
    .X(clknet_1_0__leaf_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net307 (.A(clknet_0_net307),
    .X(clknet_1_1__leaf_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net210 (.A(net210),
    .X(clknet_0_net210));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net210 (.A(clknet_0_net210),
    .X(clknet_1_0__leaf_net210));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net210 (.A(clknet_0_net210),
    .X(clknet_1_1__leaf_net210));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net187 (.A(net187),
    .X(clknet_0_net187));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net187 (.A(clknet_0_net187),
    .X(clknet_1_0__leaf_net187));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net187 (.A(clknet_0_net187),
    .X(clknet_1_1__leaf_net187));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net690 (.A(net690),
    .X(clknet_0_net690));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net690 (.A(clknet_0_net690),
    .X(clknet_1_0__leaf_net690));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net690 (.A(clknet_0_net690),
    .X(clknet_1_1__leaf_net690));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net880 (.A(net880),
    .X(clknet_0_net880));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net880 (.A(clknet_0_net880),
    .X(clknet_1_0__leaf_net880));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net880 (.A(clknet_0_net880),
    .X(clknet_1_1__leaf_net880));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net183 (.A(net183),
    .X(clknet_0_net183));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net183 (.A(clknet_0_net183),
    .X(clknet_1_0__leaf_net183));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net183 (.A(clknet_0_net183),
    .X(clknet_1_1__leaf_net183));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net689 (.A(net689),
    .X(clknet_0_net689));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net689 (.A(clknet_0_net689),
    .X(clknet_1_0__leaf_net689));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net689 (.A(clknet_0_net689),
    .X(clknet_1_1__leaf_net689));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net910 (.A(net910),
    .X(clknet_0_net910));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net910 (.A(clknet_0_net910),
    .X(clknet_1_0__leaf_net910));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net910 (.A(clknet_0_net910),
    .X(clknet_1_1__leaf_net910));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net673 (.A(net673),
    .X(clknet_0_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net673 (.A(clknet_0_net673),
    .X(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net673 (.A(clknet_0_net673),
    .X(clknet_1_1__leaf_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net224 (.A(net224),
    .X(clknet_0_net224));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net224 (.A(clknet_0_net224),
    .X(clknet_1_0__leaf_net224));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net224 (.A(clknet_0_net224),
    .X(clknet_1_1__leaf_net224));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net649 (.A(net649),
    .X(clknet_0_net649));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net649 (.A(clknet_0_net649),
    .X(clknet_1_0__leaf_net649));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net649 (.A(clknet_0_net649),
    .X(clknet_1_1__leaf_net649));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net925 (.A(net925),
    .X(clknet_0_net925));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net925 (.A(clknet_0_net925),
    .X(clknet_1_0__leaf_net925));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net925 (.A(clknet_0_net925),
    .X(clknet_1_1__leaf_net925));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net304 (.A(net304),
    .X(clknet_0_net304));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net304 (.A(clknet_0_net304),
    .X(clknet_1_0__leaf_net304));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net304 (.A(net1055),
    .X(clknet_1_1__leaf_net304));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net529 (.A(net529),
    .X(clknet_0_net529));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net529 (.A(clknet_0_net529),
    .X(clknet_1_0__leaf_net529));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net529 (.A(clknet_0_net529),
    .X(clknet_1_1__leaf_net529));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net202 (.A(net202),
    .X(clknet_0_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net202 (.A(clknet_0_net202),
    .X(clknet_1_0__leaf_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net202 (.A(clknet_0_net202),
    .X(clknet_1_1__leaf_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net922 (.A(net922),
    .X(clknet_0_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net922 (.A(clknet_0_net922),
    .X(clknet_1_0__leaf_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net922 (.A(clknet_0_net922),
    .X(clknet_1_1__leaf_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net100 (.A(net100),
    .X(clknet_0_net100));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net100 (.A(clknet_0_net100),
    .X(clknet_1_0__leaf_net100));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net100 (.A(clknet_0_net100),
    .X(clknet_1_1__leaf_net100));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net892 (.A(net892),
    .X(clknet_0_net892));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net892 (.A(clknet_0_net892),
    .X(clknet_1_0__leaf_net892));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net892 (.A(clknet_0_net892),
    .X(clknet_1_1__leaf_net892));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net672 (.A(net672),
    .X(clknet_0_net672));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net672 (.A(clknet_0_net672),
    .X(clknet_1_0__leaf_net672));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net672 (.A(clknet_0_net672),
    .X(clknet_1_1__leaf_net672));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net94 (.A(net94),
    .X(clknet_0_net94));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net94 (.A(clknet_0_net94),
    .X(clknet_1_0__leaf_net94));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net94 (.A(clknet_0_net94),
    .X(clknet_1_1__leaf_net94));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net325 (.A(net325),
    .X(clknet_0_net325));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net325 (.A(clknet_0_net325),
    .X(clknet_1_0__leaf_net325));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net325 (.A(clknet_0_net325),
    .X(clknet_1_1__leaf_net325));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net671 (.A(net671),
    .X(clknet_0_net671));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net671 (.A(clknet_0_net671),
    .X(clknet_1_0__leaf_net671));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net671 (.A(clknet_0_net671),
    .X(clknet_1_1__leaf_net671));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net88 (.A(net88),
    .X(clknet_0_net88));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net88 (.A(clknet_0_net88),
    .X(clknet_1_0__leaf_net88));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net88 (.A(clknet_0_net88),
    .X(clknet_1_1__leaf_net88));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net26),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net1034),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net1034),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net1036),
    .X(net1037));
 sky130_fd_sc_hd__mux4_1 clone5 (.A0(net976),
    .A1(net24),
    .A2(net1085),
    .A3(net982),
    .S0(net1067),
    .S1(net977),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net31),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net23),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net30),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net63),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net1042),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net63),
    .X(net1044));
 sky130_fd_sc_hd__clkbuf_4 clone12 (.A(net1046),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net28),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net1046),
    .X(net1047));
 sky130_fd_sc_hd__buf_2 rebuffer15 (.A(net1047),
    .X(net1048));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer16 (.A(net25),
    .X(net1049));
 sky130_fd_sc_hd__clkbuf_1 clone17 (.A(net23),
    .X(net1050));
 sky130_fd_sc_hd__clkbuf_4 clone18 (.A(net1052),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net31),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net969),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net1053),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(clknet_0_net304),
    .X(net1055));
 sky130_fd_sc_hd__a41o_1 clone23 (.A1(net976),
    .A2(net767),
    .A3(net18),
    .A4(net1057),
    .B1(net977),
    .X(net1056));
 sky130_fd_sc_hd__buf_4 clone24 (.A(net865),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net865),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(clknet_0_net314),
    .X(net1059));
 sky130_fd_sc_hd__clkbuf_1 clone27 (.A(net27),
    .X(net1060));
 sky130_fd_sc_hd__clkbuf_1 clone28 (.A(net21),
    .X(net1061));
 sky130_fd_sc_hd__clkbuf_1 clone29 (.A(net16),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(net1105),
    .X(net1063));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer31 (.A(net1063),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(net1064),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(net1064),
    .X(net1066));
 sky130_fd_sc_hd__clkbuf_1 clone34 (.A(net1020),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net699),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net706),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net583),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net160),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net141),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net753),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net750),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net996),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net565),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net742),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net653),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net885),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net687),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net646),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net687),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net688),
    .X(net1084));
 sky130_fd_sc_hd__buf_4 fanout1 (.A(net977),
    .X(net1068));
 sky130_fd_sc_hd__buf_12 fanout2 (.A(net980),
    .X(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in62));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in63));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in64));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(in65));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(in66));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(in67));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(in68));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(in69));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(in70));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(in71));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(in72));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(in73));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(in74));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(in75));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(in76));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(in77));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(in78));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(in79));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(in80));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(in81));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(in82));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(in83));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(in84));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(in85));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(in86));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(in87));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(in88));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(in89));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(in90));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(in91));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(in92));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(in93));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(in94));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(in95));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(in96));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(in97));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(in98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(in99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A0 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_S0 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_X (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A4 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_SCE (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_X (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_S0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_X (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A0 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A3 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A0 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_SCD (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_SCD (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_X (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_SCD (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A3 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_S0 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_Q_N (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_X (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A3 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_RESET_B (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_X (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A3 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_SCD (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_SCD (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_X (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A3 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_Q_N (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_A4 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_Q (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A0 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A0 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_SET_B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A0 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A0 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_X (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A0 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A3 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_X (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold40_A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_Q_N (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A0 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A0 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_Q (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S0 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S0 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A3 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_Q_N (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A0 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_Q (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A0 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_S0 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_X (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A3 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A3 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A3 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_Q_N (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A0 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A0 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_Q (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A0 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A3 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A3 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_S1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_X (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A0 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A4 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A2 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A2 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_RESET_B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_SCE (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A3 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_S0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_X (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A0 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A1 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A1 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A1 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A3 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A2 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A1 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A2 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A2 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A0 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_X (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A0 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A3 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A0 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A0 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_S0 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_X (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A0 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A0 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_S1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_RESET_B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_X (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A0 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A0 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_SCE (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_X (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone29_A (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_RESET_B (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_X (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A3 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_S0 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A0 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A0 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A3 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_RESET_B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_X (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A0 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A0 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A0 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_X (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A4 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A0 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A4 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A0 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_S0 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A4 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_X (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_S1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A0 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_S1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_X (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A0 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A3 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A0 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A0 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_X (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone23_A3 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A0 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A3 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S0 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A3 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_X (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_X (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A3 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_X (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_S0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_X (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_X (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone28_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_X (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone17_A (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A4 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S0 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_SCE (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_Q_N (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_Q (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A0 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A3 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A3 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_X (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A2 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A3 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A3 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A3 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_Q_N (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_Q (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A0 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_X (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_SCE (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A4 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_X (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A0 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_RESET_B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_RESET_B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_X (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_D (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_X (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_SCE (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A2 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_Q_N (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_S0 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_Q (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A0 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_S0 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A3 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A3 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A0 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_X (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_RESET_B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A3 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A3 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A3 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_Q_N (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A3 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_Q (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer16_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A0 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A3 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A2 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_X (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A0 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_RESET_B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_X (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_SCD (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_S0 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_D (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_RESET_B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_X (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net259_A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_X (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_Q (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S0 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A3 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A3 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A3 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_Q (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A0 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_Q (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone27_A (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_SCD (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A3 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A0 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A0 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_Q (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A0 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S0 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A3 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_X (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A0 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A0 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A3 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A2 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S0 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_X (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A3 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_X (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A3 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A0 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_X (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A0 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A2 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_X (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A3 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A3 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A0 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A3 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_X (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_S0 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_RESET_B (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A2 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A0 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_SCE (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_X (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A3 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A2 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A2 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_SCD (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_X (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A0 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_Q (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A0 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A3 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A0 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_D (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_RESET_B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_X (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_X (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A0 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A0 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_S0 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_S0 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A4 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_X (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A3 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_S1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_D (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_S1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A4 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A3 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_X (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net364_A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_X (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A1 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A1 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A0 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_X (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A0 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A0 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A0 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_X (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A0 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A0 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_X (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_X (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A0 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A3 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_X (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A1 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_X (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_Q_N (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_Q (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_SCE (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_X (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_S0 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A3 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_S1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A3 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_X (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_D (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A3 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_X (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A3 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_X (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A0 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A0 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S0 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A3 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_SCD (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A2 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A3 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_D (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_SCD (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_X (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A3 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A0 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A2 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A2 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_Q (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A0 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A3 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A3 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S0 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A3 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_X (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A0 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_X (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_S0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_X (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A3 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_D (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A0 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A3 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_SCD (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_X (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A3 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A0 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A3 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_S0 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_S0 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_X (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A0 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A3 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A4 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A4 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_X (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A0 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A3 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_X (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_Q (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_SCE (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A3 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S0 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A3 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_S1 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_S0 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_Q (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S1 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A1 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A3 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_Q (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A4 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A3 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A3 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_SET_B (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_Q (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A3 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A3 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A3 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A0 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_X (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_Q (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A2 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A3 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A3 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S0 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_S1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_Q (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_S1 (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_B1 (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_S0 (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A2 (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A3 (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_S1 (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A3 (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_B1 (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_Q (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A3 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A3 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S0 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A0 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A3 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A0 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_X (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_Q (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A2 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_S0 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_S0 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_S0 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S0 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_Q_N (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_S1 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A3 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A3 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_S0 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S0 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_S0 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_S0 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_S0 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S0 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S0 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A4 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S0 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A0 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A0 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A3 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A3 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A3 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A3 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_X (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S0 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S0 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_S0 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A2 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_S0 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_S1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_S0 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A0 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_X (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge848_Q (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A2 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A3 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_S0 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S1 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A0 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A3 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A0 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_S0 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A0 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_X (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_Q (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S0 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A3 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A1 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A3 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge854_Q (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A1 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A1 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_Q (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S0 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_S0 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A3 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A3 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_S0 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer11_A (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer9_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A0 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A3 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_X (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_Q (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_S1 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_S1 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S0 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S0 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge860_Q (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A2 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A3 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_Q (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S1 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A2 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A3 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_Q (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S0 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S0 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge864_Q (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A2 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_Q (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S1 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A1 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S0 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A4 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A4 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold49_A (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_Q (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S1 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S0 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A3 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_Q_N (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_S0 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S0 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A2 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_Q (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_S0 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A3 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_B1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S0 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_Q (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S0 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S1 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S1 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A2 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_S0 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S0 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_Q (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S1 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A2 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_Q (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S0 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S0 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A3 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S0 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_Q_N (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A3 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_S1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A4 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S0 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_S1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_S1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_Q (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S0 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_S0 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S0 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_S1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_B1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_Q_N (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S0 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S0 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A2 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_B1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_Q (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_B1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_S1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_Q (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A3 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S0 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A3 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_S0 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_Q (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S0 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A3 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_S0 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_S0 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_S1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_S1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_S1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net671_A (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_GCLK (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_Q (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S0 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_S0 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S1 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_Q (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A1 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S1 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S0 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_Q_N (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S0 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_S1 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_S1 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_S1 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_Q (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S0 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S1 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S1 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A3 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S1 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_A (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S0 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S1 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A4 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_Q (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_A (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_S1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S0 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_S1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_Q (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_Q_N (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_S0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_S1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_S0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_B1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_S1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_Q (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_B1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S0 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_Q_N (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S0 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_S1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_Q (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S0 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S1 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S1 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold51_A (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_Q (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S0 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_S0 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_S0 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S0 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net689_A (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_s908_GCLK (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_Q_N (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S1 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A3 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S1 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_Q (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_S0 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S0 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S0 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_S1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_S1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_S1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_Q (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S0 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A3 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_S1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_Q (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S0 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_Q (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_S0 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_SET_B (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S0 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_S1 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_s921_Q (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A3 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_S0 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A4 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_S1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_S1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_S1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A4 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold37_A (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_s922_Q (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_SET_B (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_SCE (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S1 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_B1 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net708_A (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_s924_GCLK (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A3 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_X (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_Q (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S0 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A3 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_S1 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_Q (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_S1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_s933_Q (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S0 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S0 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A3 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_S1 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_S1 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_Q (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S0 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_S1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_s938_Q (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S0 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A3 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_S1 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B1 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_s939_Q (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_S0 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S0 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_S1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_s943_Q (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S0 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A3 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_S1 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_s947_Q (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S1 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A2 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S1 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_S0 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S1 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S1 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S0 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_S0 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_S1 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_s949_Q (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_S1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_S0 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_S1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_S1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_s950_Q (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A3 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S1 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_S0 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_s954_Q (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S1 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A3 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S1 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S1 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S1 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold41_A (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_s962_Q (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A3 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_S0 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_S1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_s965_Q (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S0 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_S0 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_S1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_s966_Q (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S1 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_S1 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_S0 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_S1 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_s968_Q (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_S1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_s969_Q (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_S1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_S1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S0 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_s970_Q (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A3 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_X (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_X (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_X (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_X (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net94_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_X (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_X (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A3 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_X (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_A (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S0 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A1 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone23_A2 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A2 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A0 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A3 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_D (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A3 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A2 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A0 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A3 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A0 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A3 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_D (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A0 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A2 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout268_A (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S0 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S0 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A2 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout266_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A0 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A4 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout264_A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A3 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A0 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A4 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A0 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_A (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_S0 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A1 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_S1 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A2 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A3 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A4 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_S0 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A2 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout261_A (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_A (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_S0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A2 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A3 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A3 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A2 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_S1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_D (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_B1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A0 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A3 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A3 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_S1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_S0 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A0 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A2 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A0 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_SCD (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A2 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A3 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_S1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_S1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A0 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A0 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A0 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A2 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A3 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A0 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A0 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S0 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A0 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A3 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A2 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_S0 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_S1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_S0 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A3 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A3 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_SET_B (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_S0 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_A3 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A2 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A3 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_X (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A0 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A3 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A3 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_S0 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_D (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A3 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A0 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A3 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_S0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A3 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A0 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A0 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A2 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A2 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A2 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A3 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A3 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_S0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A2 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A3 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_S0 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A3 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A3 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A2 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A2 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A0 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A2 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A3 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_S0 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A0 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A3 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A2 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A3 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A2 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A3 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A3 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_X (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_S0 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A3 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A4 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_B1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_S1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A2 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A3 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_S0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_B1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_B1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A3 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A3 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A2 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A0 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A2 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A2 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A3 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_X (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A4 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_S0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S1 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A1 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A2 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A2 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A2 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A1 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A2 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A2 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A2 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_X (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A3 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A2 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A2 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_A3 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A2 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_X (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_B1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_A0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A2 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_S1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_S1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_X (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A3 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_X (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A3 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A2 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_X (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A0 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A2 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A3 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_X (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A3 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_X (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A2 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A2 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_A (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_X (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_X (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S0 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A0 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A3 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A0 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_X (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A0 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A3 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_X (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_SET_B (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_S0 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_S0 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A1 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_X (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A2 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A0 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A2 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A0 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A3 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A2 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_S0 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_X (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S0 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A0 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A3 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_S0 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A0 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A2 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A2 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_X (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A3 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S0 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A2 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A2 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A3 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A3 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_S0 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_S0 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_X (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S0 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_S0 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A3 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A1 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A3 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_S0 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_X (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_S0 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A0 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_S0 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A2 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer25_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone24_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_X (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_X (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A2 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A1 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_X (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_Q (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_S0 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A2 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S0 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_S0 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S0 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_S0 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S0 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_RESET_B (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A3 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A3 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A3 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A0 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_X (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold47_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_Q (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S0 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_S1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A0 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A0 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A3 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A3 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_X (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A2 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_X (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_X (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_output129_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_Q (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S0 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_Q (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A3 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_output133_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_Q (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_output134_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_Q (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S0 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_Q (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S0 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S0 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S0 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_SET_B (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_output136_A (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A3 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_X (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_output137_A (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_Q_N (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A3 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_S0 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_Q (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S0 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A3 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S0 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S0 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A3 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_output139_A (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A2 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A3 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A2 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_X (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_output140_A (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_Q (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_S0 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_output141_A (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A3 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_X (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A3 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A2 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_Q (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_output144_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_Q (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_output149_A (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A2 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_X (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_output151_A (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_Q (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S0 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S0 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S1 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_S0 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_output154_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A3 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A3 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_X (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_output155_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_Q (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_S1 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_S1 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_S1 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A2 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_output156_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A2 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_S0 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A3 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A3 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_X (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_output160_A (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A2 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_S0 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A2 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A2 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_S0 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A1 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_X (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_output162_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_Q (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A4 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A3 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A3 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_output167_A (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_X (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A4 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_output172_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_Q (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A3 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_output174_A (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_S0 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A2 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A3 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A3 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_X (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_X (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A3 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A3 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A3 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_S0 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A3 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_SCE (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A3 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_X (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A3 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A3 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S0 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_SCE (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A0 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A0 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A0 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_X (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A4 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_SCD (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_SET_B (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_X (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_S0 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_S0 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A0 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_B1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A2 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_RESET_B (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_X (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A0 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_X (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A3 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A3 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A3 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A3 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A3 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A2 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_X (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A2 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A2 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_X (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A2 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_X (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A3 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A0 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_S1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_RESET_B (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A4 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A2 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_X (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A2 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S0 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_S1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A3 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A3 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A2 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A2 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A0 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_X (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_S0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_B1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_SCD (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_X (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A3 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_S1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_SET_B (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A4 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A3 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_X (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_S0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_S0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_S1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_X (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A2 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A2 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_S0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A2 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_S0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A2 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_X (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A2 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A4 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A3 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A0 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_X (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A0 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A3 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_A3 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_X (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S0 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A0 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A4 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_S0 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A4 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A4 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A3 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_X (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A0 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_S0 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A2 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_X (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_B1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_S0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer20_A (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_X (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A1 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_B1 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_SET_B (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B1 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A2 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A1 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_X (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A0 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A3 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A2 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_S1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_S1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A3 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_X (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_S0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_SCD (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A4 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A3 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A4 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_X (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S0 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A0 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A2 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A1 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_S1 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_X (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_S1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_D (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_SCD (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_SCE (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A4 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A4 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_S1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A4 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_X (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A2 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A3 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_S0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_S1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_S0 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_S1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_X (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A2 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A2 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_X (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A4 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A3 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A2 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_S1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_X (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_B1 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A1 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A1 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A0 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout2_A (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_X (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_X (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A3 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A2 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_B1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A3 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A3 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_X (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_S0 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A3 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_X (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A3 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A3 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A3 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_S1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_S1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_X (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A3 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A3 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_A (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A3 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer30_A (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_X (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A1 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B1 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_B1 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A2 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A3 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A0 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap224_X (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A3 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire225_X (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A3 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap226_X (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_S0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_S0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_X (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A2 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_SCE (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_S0 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A3 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_S0 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_S1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_S1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_X (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S0 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_S0 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S0 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A3 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_S1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_S1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S0 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_SET_B (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_B1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_X (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A2 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A3 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_S1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_S1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A3 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold43_A (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_X (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A4 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A4 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A4 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_SCE (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S0 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A3 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S0 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A4 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_X (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_RESET_B (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A3 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_X (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A3 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_output171_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_S0 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_X (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A4 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A4 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_X (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_B1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A3 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_SCD (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_SET_B (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_B1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A3 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A4 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_X (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A0 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A4 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A0 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A3 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_S1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_A4 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_X (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A2 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A2 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A4 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A2 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_X (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S0 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_X (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A4 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A3 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A3 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_X (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A2 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A1 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A1 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A3 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S0 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_B1 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_S1 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_S0 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A1 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_X (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_SCD (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A3 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A3 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_X (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_A (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_S0 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A3 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_X (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A3 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A3 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_S0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A3 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_X (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A4 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_X (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A2 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A4 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A0 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A2 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_S1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_X (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S0 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A2 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_X (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A4 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A0 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_X (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A1 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A3 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A3 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A1 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A3 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_S0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_A4 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_X (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_SCE (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A3 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A3 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_X (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A3 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S0 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A0 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_X (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A3 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_D (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A3 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_X (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A4 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_S1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_S0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_A (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_X (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_S0 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_S0 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A4 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A2 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B1 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B1 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone34_A (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_X (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S1 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A2 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_S0 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B1 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A4 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B1 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_X (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A4 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_S0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_S0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_S0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_B1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_X (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_X (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_SCE (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_S1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A3 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_X (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A3 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A3 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A4 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A3 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_S0 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A3 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_S1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_S0 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A3 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout261_X (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A0 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A2 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout262_X (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A2 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A2 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_S1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A3 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A4 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A2 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A3 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A3 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_X (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A3 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A2 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_D (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S0 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A3 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A3 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A3 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A2 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A2 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout264_X (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_S1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_S0 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A3 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A2 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A3 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A0 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_X (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A2 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A2 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_RESET_B (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A3 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A3 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_S0 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A0 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout266_X (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A4 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A2 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A2 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A3 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A1 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A0 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A1 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_S1 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A1 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A3 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_S1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_S0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_S0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A2 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_X (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A4 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A2 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_S1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout268_X (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A2 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S0 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_S0 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A2 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A3 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A0 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_S0 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_S0 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A3 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_X (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A2 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A2 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A3 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A3 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_S0 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_B1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_S0 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s911_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge854_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge885_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_SLEEP_B (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s905_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s910_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s929_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s933_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_SLEEP_B (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_SLEEP_B (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s924_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge863_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s953_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s955_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s957_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s958_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s959_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s960_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s961_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge848_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s950_SLEEP_B (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s951_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s956_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge860_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge875_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge864_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s970_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s972_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge886_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s926_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s945_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s946_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s949_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge877_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s921_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s922_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s938_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s939_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s940_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s941_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s942_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s943_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s944_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s948_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s952_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s954_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s966_SLEEP_B (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s967_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s969_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s971_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A3 (.DIODE(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A0 (.DIODE(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S0 (.DIODE(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net887_X (.DIODE(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S1 (.DIODE(clknet_1_0__leaf_net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S0 (.DIODE(clknet_1_0__leaf_net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S0 (.DIODE(clknet_1_0__leaf_net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S0 (.DIODE(clknet_1_0__leaf_net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S1 (.DIODE(clknet_1_0__leaf_net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S0 (.DIODE(clknet_1_0__leaf_net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(clknet_1_0__leaf_net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net727_X (.DIODE(clknet_1_0__leaf_net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_B1 (.DIODE(clknet_1_1__leaf_net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_S1 (.DIODE(clknet_1_1__leaf_net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_B1 (.DIODE(clknet_1_1__leaf_net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_B1 (.DIODE(clknet_1_1__leaf_net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_S0 (.DIODE(clknet_1_1__leaf_net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_S1 (.DIODE(clknet_1_1__leaf_net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_S1 (.DIODE(clknet_1_1__leaf_net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_B1 (.DIODE(clknet_1_1__leaf_net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_S0 (.DIODE(clknet_1_1__leaf_net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net727_X (.DIODE(clknet_1_1__leaf_net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(clknet_1_0__leaf_net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A2 (.DIODE(clknet_1_0__leaf_net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(clknet_1_0__leaf_net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net382_X (.DIODE(clknet_1_0__leaf_net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net875_A (.DIODE(clknet_0_net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net875_A (.DIODE(clknet_0_net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net875_X (.DIODE(clknet_0_net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A3 (.DIODE(clknet_1_0__leaf_net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A3 (.DIODE(clknet_1_0__leaf_net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A2 (.DIODE(clknet_1_0__leaf_net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S1 (.DIODE(clknet_1_0__leaf_net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(clknet_1_0__leaf_net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net875_X (.DIODE(clknet_1_0__leaf_net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_B1 (.DIODE(clknet_1_1__leaf_net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_S1 (.DIODE(clknet_1_1__leaf_net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S1 (.DIODE(clknet_1_1__leaf_net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S1 (.DIODE(clknet_1_1__leaf_net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_S0 (.DIODE(clknet_1_1__leaf_net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A2 (.DIODE(clknet_1_1__leaf_net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net875_X (.DIODE(clknet_1_1__leaf_net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A2 (.DIODE(clknet_1_0__leaf_net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A3 (.DIODE(clknet_1_0__leaf_net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A2 (.DIODE(clknet_1_0__leaf_net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A1 (.DIODE(clknet_1_0__leaf_net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(clknet_1_0__leaf_net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net278_X (.DIODE(clknet_1_0__leaf_net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A1 (.DIODE(clknet_1_1__leaf_net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A2 (.DIODE(clknet_1_1__leaf_net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A2 (.DIODE(clknet_1_1__leaf_net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A0 (.DIODE(clknet_1_1__leaf_net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net278_X (.DIODE(clknet_1_1__leaf_net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A2 (.DIODE(clknet_1_0__leaf_net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A2 (.DIODE(clknet_1_0__leaf_net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A2 (.DIODE(clknet_1_0__leaf_net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A1 (.DIODE(clknet_1_0__leaf_net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A1 (.DIODE(clknet_1_0__leaf_net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A1 (.DIODE(clknet_1_0__leaf_net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net293_X (.DIODE(clknet_1_0__leaf_net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(clknet_1_1__leaf_net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A1 (.DIODE(clknet_1_1__leaf_net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(clknet_1_1__leaf_net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A1 (.DIODE(clknet_1_1__leaf_net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net293_X (.DIODE(clknet_1_1__leaf_net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A2 (.DIODE(clknet_1_0__leaf_net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A3 (.DIODE(clknet_1_0__leaf_net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(clknet_1_0__leaf_net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(clknet_1_0__leaf_net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net259_X (.DIODE(clknet_1_0__leaf_net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S1 (.DIODE(clknet_1_0__leaf_net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S1 (.DIODE(clknet_1_0__leaf_net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A3 (.DIODE(clknet_1_0__leaf_net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S0 (.DIODE(clknet_1_0__leaf_net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net691_X (.DIODE(clknet_1_0__leaf_net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(clknet_1_1__leaf_net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_S0 (.DIODE(clknet_1_1__leaf_net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A3 (.DIODE(clknet_1_1__leaf_net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A2 (.DIODE(clknet_1_1__leaf_net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net691_X (.DIODE(clknet_1_1__leaf_net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A2 (.DIODE(clknet_1_0__leaf_net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(clknet_1_0__leaf_net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A2 (.DIODE(clknet_1_0__leaf_net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A3 (.DIODE(clknet_1_0__leaf_net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net185_X (.DIODE(clknet_1_0__leaf_net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A0 (.DIODE(clknet_1_1__leaf_net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A0 (.DIODE(clknet_1_1__leaf_net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A0 (.DIODE(clknet_1_1__leaf_net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A0 (.DIODE(clknet_1_1__leaf_net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net185_X (.DIODE(clknet_1_1__leaf_net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A1 (.DIODE(clknet_1_0__leaf_net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A3 (.DIODE(clknet_1_0__leaf_net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net868_X (.DIODE(clknet_1_0__leaf_net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S0 (.DIODE(clknet_1_0__leaf_net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S1 (.DIODE(clknet_1_0__leaf_net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_output147_A (.DIODE(clknet_1_0__leaf_net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net911_X (.DIODE(clknet_1_0__leaf_net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S0 (.DIODE(clknet_1_1__leaf_net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A3 (.DIODE(clknet_1_1__leaf_net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(clknet_1_1__leaf_net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A3 (.DIODE(clknet_1_1__leaf_net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net911_X (.DIODE(clknet_1_1__leaf_net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net689_A (.DIODE(clknet_0_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net689_A (.DIODE(clknet_0_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net689_X (.DIODE(clknet_0_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_S1 (.DIODE(clknet_1_0__leaf_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S0 (.DIODE(clknet_1_0__leaf_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S1 (.DIODE(clknet_1_0__leaf_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A2 (.DIODE(clknet_1_0__leaf_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S0 (.DIODE(clknet_1_0__leaf_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S0 (.DIODE(clknet_1_0__leaf_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(clknet_1_0__leaf_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S1 (.DIODE(clknet_1_0__leaf_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A3 (.DIODE(clknet_1_0__leaf_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net689_X (.DIODE(clknet_1_0__leaf_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_S0 (.DIODE(clknet_1_1__leaf_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S0 (.DIODE(clknet_1_1__leaf_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S0 (.DIODE(clknet_1_1__leaf_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A3 (.DIODE(clknet_1_1__leaf_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(clknet_1_1__leaf_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S1 (.DIODE(clknet_1_1__leaf_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S0 (.DIODE(clknet_1_1__leaf_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net689_X (.DIODE(clknet_1_1__leaf_net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S0 (.DIODE(clknet_1_0__leaf_net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(clknet_1_0__leaf_net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(clknet_1_0__leaf_net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net649_X (.DIODE(clknet_1_0__leaf_net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_S1 (.DIODE(clknet_1_0__leaf_net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_S1 (.DIODE(clknet_1_0__leaf_net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_S0 (.DIODE(clknet_1_0__leaf_net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S0 (.DIODE(clknet_1_0__leaf_net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S1 (.DIODE(clknet_1_0__leaf_net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net672_X (.DIODE(clknet_1_0__leaf_net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S1 (.DIODE(clknet_1_1__leaf_net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_S1 (.DIODE(clknet_1_1__leaf_net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_S0 (.DIODE(clknet_1_1__leaf_net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S1 (.DIODE(clknet_1_1__leaf_net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_S1 (.DIODE(clknet_1_1__leaf_net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S0 (.DIODE(clknet_1_1__leaf_net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net672_X (.DIODE(clknet_1_1__leaf_net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net671_A (.DIODE(clknet_0_net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net671_A (.DIODE(clknet_0_net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net671_X (.DIODE(clknet_0_net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_S1 (.DIODE(clknet_1_0__leaf_net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S1 (.DIODE(clknet_1_0__leaf_net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S0 (.DIODE(clknet_1_0__leaf_net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S1 (.DIODE(clknet_1_0__leaf_net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net671_X (.DIODE(clknet_1_0__leaf_net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(clknet_1_1__leaf_net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S0 (.DIODE(clknet_1_1__leaf_net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S0 (.DIODE(clknet_1_1__leaf_net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S0 (.DIODE(clknet_1_1__leaf_net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net671_X (.DIODE(clknet_1_1__leaf_net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A0 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A0 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A1 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer4_X (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A3 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A2 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone5_X (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer6_X (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer8_X (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A2 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A0 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A0 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_SCE (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A0 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer10_A (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer9_X (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A0 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A2 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A2 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S0 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone12_X (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer14_A (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone12_A (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer13_X (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A3 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_S1 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A0 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A0 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A3 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone17_X (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A3 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A2 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_S0 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A2 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_RESET_B (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone18_X (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone23_A4 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A1 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A1 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A2 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A3 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A2 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone24_X (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_A (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer25_X (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A0 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A1 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A2 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A2 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A3 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone27_X (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_B1 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A0 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_SCE (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_S1 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_SCD (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone28_X (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A0 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S0 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A3 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_D (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A2 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone29_X (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer33_A (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer32_A (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer31_X (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone5_S0 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B1 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A3 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_S0 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S1 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone34_X (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_S1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold47_X (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout2_X (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone5_A2 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A3 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A2 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A3 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net817));
 sky130_fd_sc_hd__mux4_1 clone1 (.A0(net22),
    .A1(net767),
    .A2(net1000),
    .A3(net982),
    .S0(net1094),
    .S1(net1068),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net872),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net872),
    .X(net1088));
 sky130_fd_sc_hd__mux4_1 clone13 (.A0(net971),
    .A1(net150),
    .A2(net36),
    .A3(net780),
    .S0(net924),
    .S1(net959),
    .X(net1089));
 sky130_fd_sc_hd__mux4_1 clone14 (.A0(net770),
    .A1(net963),
    .A2(net1015),
    .A3(net786),
    .S0(net966),
    .S1(net970),
    .X(net1090));
 sky130_fd_sc_hd__a41o_1 clone15 (.A1(net998),
    .A2(net1001),
    .A3(net770),
    .A4(net1031),
    .B1(net1004),
    .X(net1091));
 sky130_fd_sc_hd__a41o_1 clone16 (.A1(net1014),
    .A2(net1031),
    .A3(net1005),
    .A4(net1001),
    .B1(net1110),
    .X(net1092));
 sky130_fd_sc_hd__clkbuf_1 clone19 (.A(net776),
    .X(net1093));
 sky130_fd_sc_hd__a41o_1 clone20 (.A1(net998),
    .A2(net1001),
    .A3(net770),
    .A4(net1031),
    .B1(net1004),
    .X(net1094));
 sky130_fd_sc_hd__clkbuf_1 clone21 (.A(net771),
    .X(net1095));
 sky130_fd_sc_hd__a41o_1 clone22 (.A1(net1100),
    .A2(net999),
    .A3(net1030),
    .A4(net1000),
    .B1(net1028),
    .X(net1096));
 sky130_fd_sc_hd__mux4_1 clone25 (.A0(net786),
    .A1(net56),
    .A2(net55),
    .A3(net812),
    .S0(net1032),
    .S1(net970),
    .X(net1097));
 sky130_fd_sc_hd__mux4_1 clone26 (.A0(net976),
    .A1(net24),
    .A2(net1085),
    .A3(net982),
    .S0(net1019),
    .S1(net1068),
    .X(net1098));
 sky130_fd_sc_hd__a41o_1 clone30 (.A1(net26),
    .A2(net18),
    .A3(net1000),
    .A4(net978),
    .B1(net1049),
    .X(net1099));
 sky130_fd_sc_hd__a41o_1 clone31 (.A1(net1014),
    .A2(net1031),
    .A3(net1005),
    .A4(net1001),
    .B1(net1019),
    .X(net1100));
 sky130_fd_sc_hd__clkbuf_1 clone32 (.A(net30),
    .X(net1101));
 sky130_fd_sc_hd__clkbuf_1 clone33 (.A(net31),
    .X(net1102));
 sky130_fd_sc_hd__clkbuf_1 clone35 (.A(net30),
    .X(net1103));
 sky130_fd_sc_hd__clkbuf_1 clone36 (.A(net21),
    .X(net1104));
 sky130_fd_sc_hd__clkbuf_2 rebuffer37 (.A(net986),
    .X(net1105));
 sky130_fd_sc_hd__clkbuf_1 clone38 (.A(net980),
    .X(net1106));
 sky130_fd_sc_hd__clkbuf_1 clone39 (.A(net788),
    .X(net1107));
 sky130_fd_sc_hd__clkbuf_1 clone40 (.A(net19),
    .X(net1108));
 sky130_fd_sc_hd__clkbuf_1 clone41 (.A(net27),
    .X(net1109));
 sky130_fd_sc_hd__clkbuf_1 clone42 (.A(net1111),
    .X(net1110));
 sky130_fd_sc_hd__clkbuf_1 clone43 (.A(net788),
    .X(net1111));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
