module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_0_net646;
 wire clknet_1_0__leaf_net646;
 wire clknet_1_1__leaf_net646;
 wire clknet_0_net736;
 wire clknet_1_0__leaf_net736;
 wire clknet_1_1__leaf_net736;
 wire clknet_0_net632;
 wire clknet_1_0__leaf_net632;
 wire clknet_1_1__leaf_net632;
 wire clknet_0_net735;
 wire clknet_1_0__leaf_net735;
 wire clknet_1_1__leaf_net735;
 wire clknet_0_net716;
 wire clknet_1_0__leaf_net716;
 wire clknet_1_1__leaf_net716;
 wire clknet_0_net580;
 wire clknet_1_0__leaf_net580;
 wire clknet_1_1__leaf_net580;
 wire clknet_0_net576;
 wire clknet_1_0__leaf_net576;
 wire clknet_1_1__leaf_net576;
 wire clknet_0_net577;
 wire clknet_1_0__leaf_net577;
 wire clknet_1_1__leaf_net577;
 wire clknet_0_net598;
 wire clknet_1_0__leaf_net598;
 wire clknet_1_1__leaf_net598;
 wire clknet_0_net834;
 wire clknet_1_0__leaf_net834;
 wire clknet_1_1__leaf_net834;
 wire clknet_0_net531;
 wire clknet_1_0__leaf_net531;
 wire clknet_1_1__leaf_net531;
 wire clknet_0_net702;
 wire clknet_1_0__leaf_net702;
 wire clknet_1_1__leaf_net702;
 wire clknet_0_net826;
 wire clknet_1_0__leaf_net826;
 wire clknet_1_1__leaf_net826;
 wire clknet_0_net687;
 wire clknet_1_0__leaf_net687;
 wire clknet_1_1__leaf_net687;
 wire clknet_0_net846;
 wire clknet_1_0__leaf_net846;
 wire clknet_1_1__leaf_net846;
 wire clknet_0_net501;
 wire clknet_1_0__leaf_net501;
 wire clknet_1_1__leaf_net501;
 wire clknet_0_net386;
 wire clknet_1_0__leaf_net386;
 wire clknet_1_1__leaf_net386;
 wire clknet_0_net633;
 wire clknet_1_0__leaf_net633;
 wire clknet_1_1__leaf_net633;
 wire clknet_0_net393;
 wire clknet_1_0__leaf_net393;
 wire clknet_1_1__leaf_net393;
 wire clknet_0_net389;
 wire clknet_1_0__leaf_net389;
 wire clknet_1_1__leaf_net389;
 wire clknet_0_net686;
 wire clknet_1_0__leaf_net686;
 wire clknet_1_1__leaf_net686;
 wire clknet_0_net672;
 wire clknet_1_0__leaf_net672;
 wire clknet_1_1__leaf_net672;
 wire clknet_0_net403;
 wire clknet_1_0__leaf_net403;
 wire clknet_1_1__leaf_net403;
 wire clknet_0_net831;
 wire clknet_1_0__leaf_net831;
 wire clknet_1_1__leaf_net831;
 wire clknet_0_net871;
 wire clknet_1_0__leaf_net871;
 wire clknet_1_1__leaf_net871;
 wire clknet_0_net671;
 wire clknet_1_0__leaf_net671;
 wire clknet_1_1__leaf_net671;
 wire clknet_0_net655;
 wire clknet_1_0__leaf_net655;
 wire clknet_1_1__leaf_net655;
 wire clknet_0_net299;
 wire clknet_1_0__leaf_net299;
 wire clknet_1_1__leaf_net299;
 wire clknet_0_net154;
 wire clknet_1_0__leaf_net154;
 wire clknet_1_1__leaf_net154;
 wire clknet_0_net275;
 wire clknet_1_0__leaf_net275;
 wire clknet_1_1__leaf_net275;
 wire clknet_0_net281;
 wire clknet_1_0__leaf_net281;
 wire clknet_1_1__leaf_net281;
 wire clknet_0_net280;
 wire clknet_1_0__leaf_net280;
 wire clknet_1_1__leaf_net280;
 wire clknet_0_net654;
 wire clknet_1_0__leaf_net654;
 wire clknet_1_1__leaf_net654;
 wire clknet_0_net855;
 wire clknet_1_0__leaf_net855;
 wire clknet_1_1__leaf_net855;
 wire clknet_0_net404;
 wire clknet_1_0__leaf_net404;
 wire clknet_1_1__leaf_net404;
 wire clknet_0_net859;
 wire clknet_1_0__leaf_net859;
 wire clknet_1_1__leaf_net859;
 wire clknet_0_net874;
 wire clknet_1_0__leaf_net874;
 wire clknet_1_1__leaf_net874;
 wire clknet_0_net196;
 wire clknet_1_0__leaf_net196;
 wire clknet_1_1__leaf_net196;
 wire clknet_0_net156;
 wire clknet_1_0__leaf_net156;
 wire clknet_1_1__leaf_net156;
 wire clknet_0_net155;
 wire clknet_1_0__leaf_net155;
 wire clknet_1_1__leaf_net155;
 wire clknet_0_net130;
 wire clknet_1_0__leaf_net130;
 wire clknet_1_1__leaf_net130;
 wire clknet_0_net375;
 wire clknet_1_0__leaf_net375;
 wire clknet_1_1__leaf_net375;
 wire clknet_0_net373;
 wire clknet_1_0__leaf_net373;
 wire clknet_1_1__leaf_net373;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;

 sky130_fd_sc_hd__xnor2_1 c100 (.A(net37),
    .B(net31),
    .Y(net38));
 sky130_fd_sc_hd__mux4_1 c101 (.A0(net27),
    .A1(net33),
    .A2(net22),
    .A3(net18),
    .S0(net16),
    .S1(net38),
    .X(net39));
 sky130_fd_sc_hd__a21bo_1 c102 (.A1(net31),
    .A2(net34),
    .B1_N(net37),
    .X(net40));
 sky130_fd_sc_hd__mux4_1 c103 (.A0(net23),
    .A1(net38),
    .A2(net35),
    .A3(net25),
    .S0(net40),
    .S1(net993),
    .X(net41));
 sky130_fd_sc_hd__sdfrbp_1 c104 (.CLK(clknet_leaf_7_clk),
    .D(net36),
    .RESET_B(net37),
    .SCD(net40),
    .SCE(net31),
    .Q(net43),
    .Q_N(net42));
 sky130_fd_sc_hd__xnor2_1 c105 (.A(net779),
    .B(net36),
    .Y(net44));
 sky130_fd_sc_hd__xnor2_1 c106 (.A(net31),
    .B(net19),
    .Y(net45));
 sky130_fd_sc_hd__xnor2_1 c107 (.A(net29),
    .B(net30),
    .Y(net46));
 sky130_fd_sc_hd__xnor2_1 c108 (.A(net45),
    .B(net651),
    .Y(net47));
 sky130_fd_sc_hd__dfrbp_1 c109 (.CLK(clknet_leaf_7_clk),
    .D(net40),
    .RESET_B(net31),
    .Q(net876),
    .Q_N(net48));
 sky130_fd_sc_hd__dfbbn_1 c110 (.CLK_N(clknet_leaf_8_clk),
    .D(net44),
    .RESET_B(net909),
    .SET_B(net652),
    .Q(net50),
    .Q_N(net49));
 sky130_fd_sc_hd__xnor2_1 c111 (.A(net36),
    .B(net768),
    .Y(net51));
 sky130_fd_sc_hd__xnor2_1 c112 (.A(net45),
    .B(net29),
    .Y(net52));
 sky130_fd_sc_hd__dfrbp_1 c113 (.CLK(clknet_leaf_8_clk),
    .D(net52),
    .RESET_B(net49),
    .Q(net54),
    .Q_N(net53));
 sky130_fd_sc_hd__dfrtn_1 c114 (.CLK_N(clknet_leaf_8_clk),
    .D(net51),
    .RESET_B(net44),
    .Q(net55));
 sky130_fd_sc_hd__sdfbbn_2 c115 (.CLK_N(clknet_leaf_7_clk),
    .D(net51),
    .RESET_B(net19),
    .SCD(net48),
    .SCE(net47),
    .SET_B(net31),
    .Q(net57),
    .Q_N(net56));
 sky130_fd_sc_hd__a31o_1 c116 (.A1(net949),
    .A2(net57),
    .A3(net29),
    .B1(net53),
    .X(net58));
 sky130_fd_sc_hd__dfbbn_1 c117 (.CLK_N(clknet_leaf_8_clk),
    .D(net57),
    .RESET_B(net52),
    .SET_B(net58),
    .Q(net862),
    .Q_N(net59));
 sky130_fd_sc_hd__xnor2_1 c118 (.A(net50),
    .B(net57),
    .Y(net830));
 sky130_fd_sc_hd__dfbbp_1 c119 (.CLK(clknet_leaf_8_clk),
    .D(net58),
    .RESET_B(net51),
    .SET_B(net44),
    .Q(net61),
    .Q_N(net60));
 sky130_fd_sc_hd__a21bo_1 c120 (.A1(net61),
    .A2(net59),
    .B1_N(net56),
    .X(net62));
 sky130_fd_sc_hd__sdfbbn_1 c121 (.CLK_N(clknet_leaf_8_clk),
    .D(net52),
    .RESET_B(net949),
    .SCD(net62),
    .SCE(net57),
    .SET_B(net61),
    .Q(net835),
    .Q_N(net63));
 sky130_fd_sc_hd__xnor2_1 c122 (.A(net862),
    .B(net33),
    .Y(net827));
 sky130_fd_sc_hd__mux4_1 c123 (.A0(net62),
    .A1(net827),
    .A2(net31),
    .A3(net19),
    .S0(net56),
    .S1(net60),
    .X(net64));
 sky130_fd_sc_hd__mux4_1 c124 (.A0(net47),
    .A1(net30),
    .A2(net827),
    .A3(net56),
    .S0(net64),
    .S1(net651),
    .X(net65));
 sky130_fd_sc_hd__mux4_1 c125 (.A0(net64),
    .A1(net827),
    .A2(net56),
    .A3(net31),
    .S0(net909),
    .S1(net982),
    .X(net66));
 sky130_fd_sc_hd__a21bo_2 c126 (.A1(net769),
    .A2(net766),
    .B1_N(net768),
    .X(net857));
 sky130_fd_sc_hd__xnor2_4 c127 (.A(net821),
    .B(net767),
    .Y(net67));
 sky130_fd_sc_hd__mux4_2 c128 (.A0(net768),
    .A1(net67),
    .A2(net763),
    .A3(net769),
    .S0(net907),
    .S1(net794),
    .X(net68));
 sky130_fd_sc_hd__xnor2_4 c129 (.A(net770),
    .B(net761),
    .Y(net69));
 sky130_fd_sc_hd__xnor2_4 c130 (.A(net766),
    .B(net805),
    .Y(net70));
 sky130_fd_sc_hd__a31o_4 c131 (.A1(net906),
    .A2(net821),
    .A3(net816),
    .B1(net767),
    .X(net71));
 sky130_fd_sc_hd__xnor2_2 c132 (.A(net819),
    .B(net761),
    .Y(net72));
 sky130_fd_sc_hd__xnor2_4 c133 (.A(net71),
    .B(net783),
    .Y(net73));
 sky130_fd_sc_hd__xnor2_4 c134 (.A(net73),
    .B(net907),
    .Y(net74));
 sky130_fd_sc_hd__a21bo_1 c135 (.A1(net72),
    .A2(net906),
    .B1_N(net765),
    .X(net75));
 sky130_fd_sc_hd__a21bo_2 c136 (.A1(net907),
    .A2(net75),
    .B1_N(net71),
    .X(net76));
 sky130_fd_sc_hd__a21bo_2 c137 (.A1(net75),
    .A2(net72),
    .B1_N(net69),
    .X(net77));
 sky130_fd_sc_hd__xnor2_2 c138 (.A(net763),
    .B(net74),
    .Y(net78));
 sky130_fd_sc_hd__a21bo_2 c139 (.A1(net783),
    .A2(net75),
    .B1_N(net907),
    .X(net79));
 sky130_fd_sc_hd__a41o_2 c140 (.A1(net72),
    .A2(net79),
    .A3(net906),
    .A4(net78),
    .B1(net907),
    .X(net80));
 sky130_fd_sc_hd__a21bo_2 c141 (.A1(net764),
    .A2(net76),
    .B1_N(net69),
    .X(net81));
 sky130_fd_sc_hd__a21bo_4 c142 (.A1(net81),
    .A2(net816),
    .B1_N(net820),
    .X(net82));
 sky130_fd_sc_hd__xnor2_2 c143 (.A(net82),
    .B(net81),
    .Y(net83));
 sky130_fd_sc_hd__a21bo_2 c144 (.A1(net77),
    .A2(net771),
    .B1_N(net83),
    .X(net84));
 sky130_fd_sc_hd__mux4_2 c145 (.A0(net78),
    .A1(net73),
    .A2(net764),
    .A3(net82),
    .S0(net769),
    .S1(net69),
    .X(net85));
 sky130_fd_sc_hd__mux4_2 c146 (.A0(net80),
    .A1(net85),
    .A2(net83),
    .A3(net72),
    .S0(net73),
    .S1(net82),
    .X(net86));
 sky130_fd_sc_hd__a21bo_1 c147 (.A1(net786),
    .A2(net791),
    .B1_N(net771),
    .X(net87));
 sky130_fd_sc_hd__xnor2_2 c148 (.A(net78),
    .B(net782),
    .Y(net88));
 sky130_fd_sc_hd__a21bo_1 c149 (.A1(net767),
    .A2(net84),
    .B1_N(net760),
    .X(net89));
 sky130_fd_sc_hd__xnor2_2 c150 (.A(net791),
    .B(net767),
    .Y(net90));
 sky130_fd_sc_hd__a21bo_1 c151 (.A1(net88),
    .A2(net768),
    .B1_N(net89),
    .X(net91));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net87),
    .A1(net89),
    .A2(net767),
    .A3(net69),
    .S0(net768),
    .S1(net792),
    .X(net92));
 sky130_fd_sc_hd__a21bo_1 c153 (.A1(net90),
    .A2(net87),
    .B1_N(net89),
    .X(net93));
 sky130_fd_sc_hd__xnor2_2 c154 (.A(net796),
    .B(net68),
    .Y(net94));
 sky130_fd_sc_hd__a31o_1 c155 (.A1(net68),
    .A2(net90),
    .A3(net88),
    .B1(net782),
    .X(net95));
 sky130_fd_sc_hd__a41o_1 c156 (.A1(net88),
    .A2(net79),
    .A3(net820),
    .A4(net775),
    .B1(net785),
    .X(net96));
 sky130_fd_sc_hd__xnor2_2 c157 (.A(net788),
    .B(net93),
    .Y(net97));
 sky130_fd_sc_hd__mux4_2 c158 (.A0(net93),
    .A1(net91),
    .A2(net68),
    .A3(net87),
    .S0(net789),
    .S1(net97),
    .X(net98));
 sky130_fd_sc_hd__a41o_1 c159 (.A1(net784),
    .A2(net787),
    .A3(net97),
    .A4(net780),
    .B1(net792),
    .X(net99));
 sky130_fd_sc_hd__a31o_2 c160 (.A1(net94),
    .A2(net83),
    .A3(net782),
    .B1(net787),
    .X(net100));
 sky130_fd_sc_hd__a31o_2 c161 (.A1(net790),
    .A2(net792),
    .A3(net92),
    .B1(net100),
    .X(net101));
 sky130_fd_sc_hd__mux4_2 c162 (.A0(net96),
    .A1(net101),
    .A2(net89),
    .A3(net87),
    .S0(net83),
    .S1(net99),
    .X(net102));
 sky130_fd_sc_hd__mux4_2 c163 (.A0(net778),
    .A1(net93),
    .A2(net99),
    .A3(net89),
    .S0(net98),
    .S1(net791),
    .X(net103));
 sky130_fd_sc_hd__a41o_1 c164 (.A1(net89),
    .A2(net101),
    .A3(net96),
    .A4(net887),
    .B1(net779),
    .X(net104));
 sky130_fd_sc_hd__a41o_1 c165 (.A1(net95),
    .A2(net791),
    .A3(net97),
    .A4(net104),
    .B1(net79),
    .X(net105));
 sky130_fd_sc_hd__mux4_1 c166 (.A0(net92),
    .A1(net105),
    .A2(net104),
    .A3(net90),
    .S0(net88),
    .S1(net103),
    .X(net106));
 sky130_fd_sc_hd__sdfbbp_1 c167 (.CLK(clknet_leaf_43_clk),
    .D(net100),
    .RESET_B(net106),
    .SCD(net99),
    .SCE(net782),
    .SET_B(net887),
    .Q(net108),
    .Q_N(net107));
 sky130_fd_sc_hd__a21bo_1 c168 (.A1(net771),
    .A2(net79),
    .B1_N(net0),
    .X(net109));
 sky130_fd_sc_hd__xnor2_1 c169 (.A(net91),
    .B(net782),
    .Y(net110));
 sky130_fd_sc_hd__a21bo_2 c170 (.A1(net809),
    .A2(net79),
    .B1_N(net782),
    .X(net111));
 sky130_fd_sc_hd__a21bo_2 c171 (.A1(net799),
    .A2(net109),
    .B1_N(net909),
    .X(net112));
 sky130_fd_sc_hd__xnor2_1 c172 (.A(net109),
    .B(net909),
    .Y(net113));
 sky130_fd_sc_hd__a21bo_2 c173 (.A1(net781),
    .A2(net887),
    .B1_N(net107),
    .X(net114));
 sky130_fd_sc_hd__a21bo_1 c174 (.A1(net112),
    .A2(net114),
    .B1_N(net906),
    .X(net115));
 sky130_fd_sc_hd__a21bo_1 c175 (.A1(net777),
    .A2(net111),
    .B1_N(net112),
    .X(net116));
 sky130_fd_sc_hd__a21bo_1 c176 (.A1(net99),
    .A2(net114),
    .B1_N(net110),
    .X(net117));
 sky130_fd_sc_hd__a21bo_1 c177 (.A1(net116),
    .A2(net909),
    .B1_N(net782),
    .X(net118));
 sky130_fd_sc_hd__xnor2_1 c178 (.A(net118),
    .B(net115),
    .Y(net119));
 sky130_fd_sc_hd__sdfxbp_1 c179 (.CLK(clknet_leaf_0_clk),
    .D(net110),
    .SCD(net115),
    .SCE(net119),
    .Q(net121),
    .Q_N(net120));
 sky130_fd_sc_hd__a21bo_2 c180 (.A1(net117),
    .A2(net118),
    .B1_N(net113),
    .X(net122));
 sky130_fd_sc_hd__sdfxbp_1 c181 (.CLK(clknet_leaf_0_clk),
    .D(net119),
    .SCD(net110),
    .SCE(net111),
    .Q(net123));
 sky130_fd_sc_hd__sdfxtp_1 c182 (.CLK(clknet_leaf_43_clk),
    .D(net965),
    .SCD(net119),
    .SCE(net776),
    .Q(net124));
 sky130_fd_sc_hd__sdfxtp_1 c183 (.CLK(clknet_leaf_0_clk),
    .D(net113),
    .SCD(net122),
    .SCE(net952),
    .Q(net125));
 sky130_fd_sc_hd__mux4_1 c184 (.A0(net952),
    .A1(net887),
    .A2(net118),
    .A3(net812),
    .S0(net109),
    .S1(net122),
    .X(net126));
 sky130_fd_sc_hd__sdfxtp_1 c185 (.CLK(clknet_leaf_43_clk),
    .D(net111),
    .SCD(net122),
    .SCE(net115),
    .Q(net127));
 sky130_fd_sc_hd__mux4_1 c186 (.A0(net97),
    .A1(net112),
    .A2(net760),
    .A3(net92),
    .S0(net118),
    .S1(net900),
    .X(net128));
 sky130_fd_sc_hd__mux4_1 c187 (.A0(net79),
    .A1(net109),
    .A2(net112),
    .A3(net906),
    .S0(net122),
    .S1(net900),
    .X(net129));
 sky130_fd_sc_hd__mux4_1 c188 (.A0(net128),
    .A1(net127),
    .A2(net797),
    .A3(net782),
    .S0(net900),
    .S1(clknet_1_0__leaf_net859),
    .X(net130));
 sky130_fd_sc_hd__sdfbbn_1 c189 (.CLK_N(clknet_leaf_5_clk),
    .D(net125),
    .RESET_B(net17),
    .SCD(net77),
    .SCE(net897),
    .SET_B(net122),
    .Q(net131));
 sky130_fd_sc_hd__a21bo_1 c190 (.A1(net1),
    .A2(net108),
    .B1_N(net13),
    .X(net132));
 sky130_fd_sc_hd__a21bo_1 c191 (.A1(net818),
    .A2(net77),
    .B1_N(net808),
    .X(net133));
 sky130_fd_sc_hd__a21bo_1 c192 (.A1(net90),
    .A2(net907),
    .B1_N(net104),
    .X(net134));
 sky130_fd_sc_hd__a21bo_1 c193 (.A1(net131),
    .A2(net17),
    .B1_N(net21),
    .X(net135));
 sky130_fd_sc_hd__a21bo_1 c194 (.A1(net18),
    .A2(net21),
    .B1_N(net792),
    .X(net136));
 sky130_fd_sc_hd__xnor2_1 c195 (.A(net134),
    .B(net136),
    .Y(net137));
 sky130_fd_sc_hd__a21bo_1 c196 (.A1(net104),
    .A2(net812),
    .B1_N(net135),
    .X(net138));
 sky130_fd_sc_hd__a21bo_1 c197 (.A1(net17),
    .A2(net804),
    .B1_N(net884),
    .X(net139));
 sky130_fd_sc_hd__a21bo_1 c198 (.A1(net808),
    .A2(net108),
    .B1_N(net900),
    .X(net140));
 sky130_fd_sc_hd__mux4_1 c199 (.A0(net20),
    .A1(net804),
    .A2(net21),
    .A3(net12),
    .S0(net135),
    .S1(net898),
    .X(net141));
 sky130_fd_sc_hd__sdfbbn_2 c200 (.CLK_N(clknet_leaf_5_clk),
    .D(net137),
    .RESET_B(net134),
    .SCD(net1),
    .SCE(net125),
    .SET_B(net898),
    .Q(net143),
    .Q_N(net142));
 sky130_fd_sc_hd__sdfbbp_1 c201 (.CLK(clknet_leaf_6_clk),
    .D(net139),
    .RESET_B(net760),
    .SCD(net898),
    .SCE(net141),
    .SET_B(net6),
    .Q(net145),
    .Q_N(net144));
 sky130_fd_sc_hd__mux4_1 c202 (.A0(net782),
    .A1(net787),
    .A2(net122),
    .A3(net901),
    .S0(net884),
    .S1(net142),
    .X(net146));
 sky130_fd_sc_hd__sdfbbn_1 c203 (.CLK_N(clknet_leaf_5_clk),
    .D(net115),
    .RESET_B(net6),
    .SCD(net898),
    .SCE(net143),
    .SET_B(net122),
    .Q(net148),
    .Q_N(net147));
 sky130_fd_sc_hd__a31o_1 c204 (.A1(net812),
    .A2(net148),
    .A3(net142),
    .B1(net898),
    .X(net149));
 sky130_fd_sc_hd__dfbbn_1 c205 (.CLK_N(clknet_leaf_5_clk),
    .D(net149),
    .RESET_B(net139),
    .SET_B(net996),
    .Q(net151),
    .Q_N(net150));
 sky130_fd_sc_hd__mux4_1 c206 (.A0(net148),
    .A1(net143),
    .A2(net898),
    .A3(net884),
    .S0(net139),
    .S1(net808),
    .X(net152));
 sky130_fd_sc_hd__mux4_1 c207 (.A0(net122),
    .A1(net901),
    .A2(net145),
    .A3(net137),
    .S0(net148),
    .S1(clknet_1_0__leaf_net655),
    .X(net153));
 sky130_fd_sc_hd__mux4_1 c208 (.A0(net133),
    .A1(net132),
    .A2(net147),
    .A3(clknet_1_0__leaf_net654),
    .S0(clknet_1_0__leaf_net655),
    .S1(net657),
    .X(net154));
 sky130_fd_sc_hd__mux4_1 c209 (.A0(net6),
    .A1(net898),
    .A2(net121),
    .A3(net147),
    .S0(clknet_1_0__leaf_net859),
    .S1(net656),
    .X(net155));
 sky130_fd_sc_hd__a21bo_1 c210 (.A1(net820),
    .A2(net34),
    .B1_N(clknet_1_0__leaf_net859),
    .X(net156));
 sky130_fd_sc_hd__xnor2_1 c211 (.A(net34),
    .B(net11),
    .Y(net157));
 sky130_fd_sc_hd__dfbbn_1 c212 (.CLK_N(clknet_leaf_7_clk),
    .D(net38),
    .RESET_B(net149),
    .SET_B(net652),
    .Q(net159),
    .Q_N(net158));
 sky130_fd_sc_hd__a21bo_1 c213 (.A1(net141),
    .A2(net159),
    .B1_N(net92),
    .X(net160));
 sky130_fd_sc_hd__a31o_2 c214 (.A1(net797),
    .A2(net909),
    .A3(net142),
    .B1(net102),
    .X(net161));
 sky130_fd_sc_hd__xnor2_1 c215 (.A(net92),
    .B(net12),
    .Y(net162));
 sky130_fd_sc_hd__dfbbp_1 c216 (.CLK(clknet_leaf_6_clk),
    .D(clknet_1_1__leaf_net156),
    .RESET_B(net161),
    .SET_B(net948),
    .Q(net164),
    .Q_N(net163));
 sky130_fd_sc_hd__sdfrbp_1 c217 (.CLK(clknet_leaf_6_clk),
    .D(clknet_1_0__leaf_net156),
    .RESET_B(net945),
    .SCD(net92),
    .SCE(net161),
    .Q(net166),
    .Q_N(net165));
 sky130_fd_sc_hd__a31o_2 c218 (.A1(net143),
    .A2(net18),
    .A3(net111),
    .B1(net160),
    .X(net167));
 sky130_fd_sc_hd__sdfxbp_1 c219 (.CLK(clknet_leaf_6_clk),
    .D(net167),
    .SCD(net18),
    .SCE(net161),
    .Q(net852),
    .Q_N(net168));
 sky130_fd_sc_hd__mux4_2 c220 (.A0(net134),
    .A1(net35),
    .A2(net92),
    .A3(net142),
    .S0(net43),
    .S1(net161),
    .X(net169));
 sky130_fd_sc_hd__sdfxbp_1 c221 (.CLK(clknet_leaf_6_clk),
    .D(net955),
    .SCD(net169),
    .SCE(net162),
    .Q(net171),
    .Q_N(net170));
 sky130_fd_sc_hd__a41o_1 c222 (.A1(net162),
    .A2(net760),
    .A3(net820),
    .A4(net170),
    .B1(net168),
    .X(net172));
 sky130_fd_sc_hd__sdfxtp_1 c223 (.CLK(clknet_leaf_6_clk),
    .D(net954),
    .SCD(net172),
    .SCE(net169),
    .Q(net173));
 sky130_fd_sc_hd__xnor2_1 c224 (.A(net161),
    .B(net898),
    .Y(net174));
 sky130_fd_sc_hd__a21bo_1 c225 (.A1(net172),
    .A2(net174),
    .B1_N(net143),
    .X(net175));
 sky130_fd_sc_hd__a21bo_2 c226 (.A1(net173),
    .A2(net165),
    .B1_N(net144),
    .X(net850));
 sky130_fd_sc_hd__a21bo_1 c227 (.A1(net11),
    .A2(net173),
    .B1_N(net850),
    .X(net176));
 sky130_fd_sc_hd__mux4_1 c228 (.A0(net43),
    .A1(net149),
    .A2(net174),
    .A3(net850),
    .S0(net175),
    .S1(net176),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 c229 (.A0(net174),
    .A1(net167),
    .A2(net175),
    .A3(net158),
    .S0(net7),
    .S1(net659),
    .X(net178));
 sky130_fd_sc_hd__mux4_1 c230 (.A0(net176),
    .A1(net850),
    .A2(net787),
    .A3(net28),
    .S0(net175),
    .S1(net869),
    .X(net179));
 sky130_fd_sc_hd__a21bo_1 c231 (.A1(net898),
    .A2(net54),
    .B1_N(net652),
    .X(net853));
 sky130_fd_sc_hd__a31o_1 c232 (.A1(net787),
    .A2(net768),
    .A3(net57),
    .B1(clknet_1_1__leaf_net859),
    .X(net180));
 sky130_fd_sc_hd__a41o_1 c233 (.A1(net159),
    .A2(net63),
    .A3(net807),
    .A4(net56),
    .B1(net853),
    .X(net181));
 sky130_fd_sc_hd__a21bo_1 c234 (.A1(net145),
    .A2(net789),
    .B1_N(net22),
    .X(net182));
 sky130_fd_sc_hd__a41o_1 c235 (.A1(net760),
    .A2(net182),
    .A3(net158),
    .A4(net898),
    .B1(net652),
    .X(net183));
 sky130_fd_sc_hd__a21bo_1 c236 (.A1(net182),
    .A2(net853),
    .B1_N(net907),
    .X(net184));
 sky130_fd_sc_hd__a31o_2 c237 (.A1(net183),
    .A2(net876),
    .A3(net768),
    .B1(net182),
    .X(net185));
 sky130_fd_sc_hd__sdfxtp_1 c238 (.CLK(clknet_leaf_7_clk),
    .D(net157),
    .SCD(net185),
    .SCE(net787),
    .Q(net186));
 sky130_fd_sc_hd__a41o_1 c239 (.A1(net768),
    .A2(net22),
    .A3(net182),
    .A4(net56),
    .B1(net186),
    .X(net187));
 sky130_fd_sc_hd__sdfbbn_1 c240 (.CLK_N(clknet_leaf_9_clk),
    .D(net46),
    .RESET_B(net145),
    .SCD(net183),
    .SCE(net185),
    .SET_B(net660),
    .Q(net841),
    .Q_N(net188));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(net181),
    .A1(net187),
    .A2(net183),
    .A3(net188),
    .S0(net167),
    .S1(net185),
    .X(net189));
 sky130_fd_sc_hd__sdfbbp_1 c242 (.CLK(clknet_leaf_9_clk),
    .D(net184),
    .RESET_B(net46),
    .SCD(net182),
    .SCE(net807),
    .SET_B(net140),
    .Q(net863));
 sky130_fd_sc_hd__a21bo_1 c243 (.A1(net185),
    .A2(net187),
    .B1_N(net163),
    .X(net190));
 sky130_fd_sc_hd__mux4_1 c244 (.A0(net180),
    .A1(net185),
    .A2(net168),
    .A3(net182),
    .S0(net59),
    .S1(clknet_1_1__leaf_net859),
    .X(net874));
 sky130_fd_sc_hd__sdfbbn_1 c245 (.CLK_N(clknet_leaf_9_clk),
    .D(net22),
    .RESET_B(clknet_1_0__leaf_net874),
    .SCD(net190),
    .SCE(net167),
    .SET_B(net660),
    .Q(net192),
    .Q_N(net191));
 sky130_fd_sc_hd__mux4_1 c246 (.A0(net54),
    .A1(net192),
    .A2(net187),
    .A3(net853),
    .S0(net188),
    .S1(net869),
    .X(net193));
 sky130_fd_sc_hd__mux4_2 c247 (.A0(net164),
    .A1(net193),
    .A2(net852),
    .A3(net190),
    .S0(net22),
    .S1(net185),
    .X(net833));
 sky130_fd_sc_hd__sdfbbn_1 c248 (.CLK_N(clknet_leaf_10_clk),
    .D(net972),
    .RESET_B(net193),
    .SCD(net144),
    .SCE(net157),
    .SET_B(net833),
    .Q(net195),
    .Q_N(net194));
 sky130_fd_sc_hd__a41o_1 c249 (.A1(net195),
    .A2(net164),
    .A3(clknet_1_0__leaf_net874),
    .A4(net190),
    .B1(net185),
    .X(net196));
 sky130_fd_sc_hd__a31o_1 c250 (.A1(net187),
    .A2(net190),
    .A3(net191),
    .B1(net194),
    .X(net836));
 sky130_fd_sc_hd__mux4_1 c251 (.A0(net175),
    .A1(clknet_1_0__leaf_net196),
    .A2(net195),
    .A3(net833),
    .S0(net188),
    .S1(net867),
    .X(net197));
 sky130_fd_sc_hd__xnor2_2 c252 (.A(net769),
    .B(net773),
    .Y(net198));
 sky130_fd_sc_hd__xnor2_4 c253 (.A(net86),
    .B(net74),
    .Y(net199));
 sky130_fd_sc_hd__xnor2_4 c254 (.A(net906),
    .B(net893),
    .Y(net200));
 sky130_fd_sc_hd__xnor2_4 c255 (.A(net76),
    .B(net816),
    .Y(net201));
 sky130_fd_sc_hd__xnor2_4 c256 (.A(net893),
    .B(net914),
    .Y(net202));
 sky130_fd_sc_hd__xnor2_4 c257 (.A(net202),
    .B(net200),
    .Y(net203));
 sky130_fd_sc_hd__a21bo_4 c258 (.A1(net816),
    .A2(net200),
    .B1_N(net203),
    .X(net204));
 sky130_fd_sc_hd__a21bo_2 c259 (.A1(net201),
    .A2(net204),
    .B1_N(net890),
    .X(net205));
 sky130_fd_sc_hd__a31o_2 c260 (.A1(net74),
    .A2(net941),
    .A3(net769),
    .B1(net890),
    .X(net206));
 sky130_fd_sc_hd__xnor2_4 c261 (.A(net773),
    .B(net67),
    .Y(net207));
 sky130_fd_sc_hd__a21bo_1 c262 (.A1(net766),
    .A2(net207),
    .B1_N(net204),
    .X(net208));
 sky130_fd_sc_hd__a41o_1 c263 (.A1(net941),
    .A2(net201),
    .A3(net893),
    .A4(net76),
    .B1(net915),
    .X(net209));
 sky130_fd_sc_hd__xnor2_4 c264 (.A(net794),
    .B(net205),
    .Y(net210));
 sky130_fd_sc_hd__mux4_2 c265 (.A0(net204),
    .A1(net915),
    .A2(net209),
    .A3(net819),
    .S0(net208),
    .S1(net942),
    .X(net211));
 sky130_fd_sc_hd__a21bo_1 c266 (.A1(net210),
    .A2(net80),
    .B1_N(net207),
    .X(net212));
 sky130_fd_sc_hd__a21bo_1 c267 (.A1(net207),
    .A2(net200),
    .B1_N(net204),
    .X(net213));
 sky130_fd_sc_hd__mux4_2 c268 (.A0(net209),
    .A1(net201),
    .A2(net212),
    .A3(net206),
    .S0(net207),
    .S1(net893),
    .X(net214));
 sky130_fd_sc_hd__sdfxtp_4 c269 (.CLK(clknet_leaf_40_clk),
    .D(net208),
    .SCD(net201),
    .SCE(net214),
    .Q(net215));
 sky130_fd_sc_hd__a21bo_1 c270 (.A1(net67),
    .A2(net213),
    .B1_N(net885),
    .X(net216));
 sky130_fd_sc_hd__mux4_2 c271 (.A0(net216),
    .A1(net215),
    .A2(net213),
    .A3(net201),
    .S0(net896),
    .S1(net207),
    .X(net217));
 sky130_fd_sc_hd__mux4_1 c272 (.A0(net205),
    .A1(net910),
    .A2(net771),
    .A3(net214),
    .S0(net939),
    .S1(net885),
    .X(net218));
 sky130_fd_sc_hd__xnor2_4 c273 (.A(net938),
    .B(net893),
    .Y(net219));
 sky130_fd_sc_hd__xnor2_4 c274 (.A(net771),
    .B(net887),
    .Y(net220));
 sky130_fd_sc_hd__xnor2_2 c275 (.A(net94),
    .B(net100),
    .Y(net221));
 sky130_fd_sc_hd__xnor2_2 c276 (.A(net775),
    .B(net780),
    .Y(net222));
 sky130_fd_sc_hd__xnor2_2 c277 (.A(net220),
    .B(net219),
    .Y(net223));
 sky130_fd_sc_hd__xnor2_4 c278 (.A(net940),
    .B(net81),
    .Y(net224));
 sky130_fd_sc_hd__xnor2_1 c279 (.A(net96),
    .B(net101),
    .Y(net225));
 sky130_fd_sc_hd__mux4_2 c280 (.A0(net212),
    .A1(net938),
    .A2(net108),
    .A3(net202),
    .S0(net219),
    .S1(net220),
    .X(net226));
 sky130_fd_sc_hd__dfrtp_4 c281 (.CLK(clknet_leaf_42_clk),
    .D(net222),
    .RESET_B(net226),
    .Q(net227));
 sky130_fd_sc_hd__a21bo_4 c282 (.A1(net200),
    .A2(net212),
    .B1_N(net220),
    .X(net228));
 sky130_fd_sc_hd__dfbbn_1 c283 (.CLK_N(clknet_leaf_42_clk),
    .D(net106),
    .RESET_B(net98),
    .SET_B(net226),
    .Q(net230),
    .Q_N(net229));
 sky130_fd_sc_hd__xnor2_1 c284 (.A(net223),
    .B(net792),
    .Y(net231));
 sky130_fd_sc_hd__a21bo_2 c285 (.A1(net222),
    .A2(net96),
    .B1_N(net224),
    .X(net232));
 sky130_fd_sc_hd__a21bo_4 c286 (.A1(net219),
    .A2(net223),
    .B1_N(net229),
    .X(net233));
 sky130_fd_sc_hd__dfrtp_4 c287 (.CLK(clknet_leaf_37_clk),
    .D(net231),
    .RESET_B(net232),
    .Q(net234));
 sky130_fd_sc_hd__sdfbbp_1 c288 (.CLK(clknet_leaf_42_clk),
    .D(net226),
    .RESET_B(net228),
    .SCD(net223),
    .SCE(net198),
    .SET_B(net893),
    .Q(net236),
    .Q_N(net235));
 sky130_fd_sc_hd__xnor2_1 c289 (.A(net234),
    .B(net235),
    .Y(net237));
 sky130_fd_sc_hd__a41o_4 c290 (.A1(net236),
    .A2(net219),
    .A3(net232),
    .A4(net221),
    .B1(net885),
    .X(net825));
 sky130_fd_sc_hd__sdfbbn_2 c291 (.CLK_N(clknet_leaf_1_clk),
    .D(net227),
    .RESET_B(net233),
    .SCD(net226),
    .SCE(net237),
    .SET_B(net825),
    .Q(net239),
    .Q_N(net238));
 sky130_fd_sc_hd__mux4_2 c292 (.A0(net237),
    .A1(net239),
    .A2(net775),
    .A3(net234),
    .S0(net225),
    .S1(net779),
    .X(net240));
 sky130_fd_sc_hd__mux4_2 c293 (.A0(net225),
    .A1(net816),
    .A2(net220),
    .A3(net240),
    .S0(net222),
    .S1(net238),
    .X(net832));
 sky130_fd_sc_hd__xnor2_2 c294 (.A(net240),
    .B(net770),
    .Y(net241));
 sky130_fd_sc_hd__dfbbn_1 c295 (.CLK_N(clknet_leaf_1_clk),
    .D(net241),
    .RESET_B(net228),
    .SET_B(net893),
    .Q(net242));
 sky130_fd_sc_hd__a21bo_1 c296 (.A1(net774),
    .A2(net103),
    .B1_N(net885),
    .X(net243));
 sky130_fd_sc_hd__xnor2_2 c297 (.A(net114),
    .B(net112),
    .Y(net244));
 sky130_fd_sc_hd__a21bo_1 c298 (.A1(net221),
    .A2(net779),
    .B1_N(net885),
    .X(net245));
 sky130_fd_sc_hd__a41o_1 c299 (.A1(net242),
    .A2(net243),
    .A3(net789),
    .A4(net234),
    .B1(net241),
    .X(net246));
 sky130_fd_sc_hd__sdfbbn_1 c300 (.CLK_N(clknet_leaf_0_clk),
    .D(net243),
    .RESET_B(net246),
    .SCD(net120),
    .SCE(net911),
    .SET_B(net234),
    .Q(net247));
 sky130_fd_sc_hd__dfbbp_1 c301 (.CLK(clknet_leaf_1_clk),
    .D(net246),
    .RESET_B(net103),
    .SET_B(net832),
    .Q(net248));
 sky130_fd_sc_hd__a21bo_2 c302 (.A1(net245),
    .A2(net114),
    .B1_N(net103),
    .X(net249));
 sky130_fd_sc_hd__xnor2_1 c303 (.A(net776),
    .B(net221),
    .Y(net250));
 sky130_fd_sc_hd__a21bo_1 c304 (.A1(net247),
    .A2(net244),
    .B1_N(net771),
    .X(net251));
 sky130_fd_sc_hd__sdfxbp_1 c305 (.CLK(clknet_leaf_1_clk),
    .D(net103),
    .SCD(net249),
    .SCE(net238),
    .Q(net252));
 sky130_fd_sc_hd__sdfxbp_1 c306 (.CLK(clknet_leaf_2_clk),
    .D(net251),
    .SCD(net249),
    .SCE(net215),
    .Q(net254),
    .Q_N(net253));
 sky130_fd_sc_hd__sdfbbp_1 c307 (.CLK(clknet_leaf_1_clk),
    .D(net250),
    .RESET_B(net251),
    .SCD(net241),
    .SCE(net893),
    .SET_B(net112),
    .Q(net256),
    .Q_N(net255));
 sky130_fd_sc_hd__a41o_1 c308 (.A1(net93),
    .A2(net800),
    .A3(net224),
    .A4(net77),
    .B1(net893),
    .X(net257));
 sky130_fd_sc_hd__sdfbbn_1 c309 (.CLK_N(clknet_leaf_1_clk),
    .D(net252),
    .RESET_B(net251),
    .SCD(net257),
    .SCE(net244),
    .SET_B(net241),
    .Q(net258));
 sky130_fd_sc_hd__sdfbbn_1 c310 (.CLK_N(clknet_leaf_1_clk),
    .D(net256),
    .RESET_B(net832),
    .SCD(net244),
    .SCE(net246),
    .SET_B(clknet_1_0__leaf_net859),
    .Q(net260),
    .Q_N(net259));
 sky130_fd_sc_hd__mux4_1 c311 (.A0(net248),
    .A1(net100),
    .A2(net259),
    .A3(net249),
    .S0(net246),
    .S1(net257),
    .X(net261));
 sky130_fd_sc_hd__sdfbbp_1 c312 (.CLK(clknet_leaf_1_clk),
    .D(net257),
    .RESET_B(clknet_1_0__leaf_net130),
    .SCD(net249),
    .SCE(net103),
    .SET_B(net663),
    .Q(net263),
    .Q_N(net262));
 sky130_fd_sc_hd__a21bo_1 c313 (.A1(net258),
    .A2(net260),
    .B1_N(net257),
    .X(net264));
 sky130_fd_sc_hd__mux4_2 c314 (.A0(net257),
    .A1(net264),
    .A2(net259),
    .A3(net215),
    .S0(net262),
    .S1(net255),
    .X(net265));
 sky130_fd_sc_hd__a21bo_1 c315 (.A1(net244),
    .A2(net803),
    .B1_N(net135),
    .X(net266));
 sky130_fd_sc_hd__sdfxtp_1 c316 (.CLK(clknet_leaf_4_clk),
    .D(clknet_1_1__leaf_net155),
    .SCD(net13),
    .SCE(net233),
    .Q(net267));
 sky130_fd_sc_hd__a21bo_1 c317 (.A1(net946),
    .A2(net243),
    .B1_N(net207),
    .X(net268));
 sky130_fd_sc_hd__mux4_1 c318 (.A0(net268),
    .A1(net239),
    .A2(net825),
    .A3(net253),
    .S0(clknet_1_0__leaf_net654),
    .S1(clknet_1_0__leaf_net655),
    .X(net269));
 sky130_fd_sc_hd__sdfxtp_1 c319 (.CLK(clknet_leaf_0_clk),
    .D(net268),
    .SCD(net77),
    .SCE(net893),
    .Q(net270));
 sky130_fd_sc_hd__a21bo_1 c320 (.A1(net267),
    .A2(net909),
    .B1_N(net657),
    .X(net271));
 sky130_fd_sc_hd__sdfrtn_1 c321 (.CLK_N(clknet_leaf_4_clk),
    .D(net991),
    .RESET_B(net268),
    .SCD(net102),
    .SCE(net804),
    .Q(net272));
 sky130_fd_sc_hd__a21bo_1 c322 (.A1(net1007),
    .A2(net272),
    .B1_N(net120),
    .X(net273));
 sky130_fd_sc_hd__a21bo_2 c323 (.A1(net273),
    .A2(net215),
    .B1_N(net238),
    .X(net274));
 sky130_fd_sc_hd__sdfxtp_1 c324 (.CLK(clknet_leaf_0_clk),
    .D(net272),
    .SCD(net244),
    .SCE(net268),
    .Q(net845));
 sky130_fd_sc_hd__a41o_1 c325 (.A1(net902),
    .A2(clknet_1_0__leaf_net154),
    .A3(net274),
    .A4(net885),
    .B1(net77),
    .X(net275));
 sky130_fd_sc_hd__a41o_1 c326 (.A1(net273),
    .A2(net271),
    .A3(net907),
    .A4(net272),
    .B1(net902),
    .X(net276));
 sky130_fd_sc_hd__a21bo_1 c327 (.A1(net270),
    .A2(net207),
    .B1_N(net271),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(net804),
    .A1(net249),
    .A2(net273),
    .A3(clknet_1_0__leaf_net275),
    .S0(net902),
    .S1(net277),
    .X(net278));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net277),
    .A1(clknet_1_0__leaf_net275),
    .A2(net265),
    .A3(clknet_1_0__leaf_net155),
    .S0(net664),
    .S1(net666),
    .X(net279));
 sky130_fd_sc_hd__mux4_1 c330 (.A0(clknet_1_0__leaf_net275),
    .A1(net761),
    .A2(net273),
    .A3(net239),
    .S0(net902),
    .S1(net656),
    .X(net280));
 sky130_fd_sc_hd__a41o_1 c331 (.A1(clknet_1_1__leaf_net275),
    .A2(net902),
    .A3(net7),
    .A4(net665),
    .B1(net667),
    .X(net281));
 sky130_fd_sc_hd__mux4_1 c332 (.A0(net274),
    .A1(net243),
    .A2(net21),
    .A3(net902),
    .S0(net664),
    .S1(net666),
    .X(net282));
 sky130_fd_sc_hd__sdfrtp_1 c333 (.CLK(clknet_leaf_3_clk),
    .D(net282),
    .RESET_B(net272),
    .SCD(net902),
    .SCE(net992),
    .Q(net283));
 sky130_fd_sc_hd__mux4_1 c334 (.A0(clknet_1_0__leaf_net280),
    .A1(net268),
    .A2(net271),
    .A3(net274),
    .S0(net902),
    .S1(net657),
    .X(net284));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(clknet_1_1__leaf_net280),
    .A1(net283),
    .A2(net802),
    .A3(net265),
    .S0(net228),
    .S1(clknet_1_1__leaf_net275),
    .X(net285));
 sky130_fd_sc_hd__a21bo_1 c336 (.A1(net239),
    .A2(net276),
    .B1_N(net875),
    .X(net286));
 sky130_fd_sc_hd__a21bo_2 c337 (.A1(net35),
    .A2(net107),
    .B1_N(net902),
    .X(net287));
 sky130_fd_sc_hd__a21bo_1 c338 (.A1(net132),
    .A2(net286),
    .B1_N(net902),
    .X(net288));
 sky130_fd_sc_hd__a21bo_2 c339 (.A1(net276),
    .A2(net7),
    .B1_N(net897),
    .X(net289));
 sky130_fd_sc_hd__a21bo_1 c340 (.A1(net160),
    .A2(net903),
    .B1_N(net163),
    .X(net290));
 sky130_fd_sc_hd__xnor2_2 c341 (.A(net207),
    .B(net287),
    .Y(net291));
 sky130_fd_sc_hd__dfbbn_1 c342 (.CLK_N(clknet_leaf_13_clk),
    .D(net254),
    .RESET_B(net290),
    .SET_B(net897),
    .Q(net293),
    .Q_N(net292));
 sky130_fd_sc_hd__mux4_1 c343 (.A0(net135),
    .A1(net27),
    .A2(net224),
    .A3(net290),
    .S0(net7),
    .S1(net903),
    .X(net294));
 sky130_fd_sc_hd__a21bo_1 c344 (.A1(net293),
    .A2(net289),
    .B1_N(net905),
    .X(net872));
 sky130_fd_sc_hd__a21bo_1 c345 (.A1(net286),
    .A2(net135),
    .B1_N(net289),
    .X(net295));
 sky130_fd_sc_hd__dfbbn_1 c346 (.CLK_N(clknet_leaf_13_clk),
    .D(net7),
    .RESET_B(net291),
    .SET_B(net290),
    .Q(net297),
    .Q_N(net296));
 sky130_fd_sc_hd__mux4_2 c347 (.A0(net108),
    .A1(net909),
    .A2(net27),
    .A3(net884),
    .S0(net287),
    .S1(net670),
    .X(net298));
 sky130_fd_sc_hd__mux4_1 c348 (.A0(net288),
    .A1(net174),
    .A2(net132),
    .A3(net903),
    .S0(net27),
    .S1(clknet_1_0__leaf_net655),
    .X(net299));
 sky130_fd_sc_hd__xnor2_1 c349 (.A(net803),
    .B(net832),
    .Y(net300));
 sky130_fd_sc_hd__a21bo_1 c350 (.A1(net295),
    .A2(net872),
    .B1_N(net660),
    .X(net838));
 sky130_fd_sc_hd__a21bo_1 c351 (.A1(net838),
    .A2(net803),
    .B1_N(net670),
    .X(net301));
 sky130_fd_sc_hd__a31o_4 c352 (.A1(net121),
    .A2(net903),
    .A3(net286),
    .B1(net107),
    .X(net822));
 sky130_fd_sc_hd__mux4_1 c353 (.A0(net301),
    .A1(net287),
    .A2(net838),
    .A3(net292),
    .S0(net884),
    .S1(net998),
    .X(net302));
 sky130_fd_sc_hd__sdfbbn_1 c354 (.CLK_N(clknet_leaf_14_clk),
    .D(net290),
    .RESET_B(net27),
    .SCD(net983),
    .SCE(net903),
    .SET_B(net825),
    .Q(net304),
    .Q_N(net303));
 sky130_fd_sc_hd__mux4_1 c355 (.A0(net304),
    .A1(net301),
    .A2(net822),
    .A3(net289),
    .S0(net238),
    .S1(net658),
    .X(net305));
 sky130_fd_sc_hd__a21bo_1 c356 (.A1(net295),
    .A2(net659),
    .B1_N(clknet_1_0__leaf_net672),
    .X(net831));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net789),
    .A1(net822),
    .A2(net833),
    .A3(net838),
    .S0(clknet_1_0__leaf_net831),
    .S1(net867),
    .X(net871));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(clknet_1_1__leaf_net871),
    .A1(clknet_1_1__leaf_net196),
    .A2(net830),
    .A3(net872),
    .S0(net867),
    .S1(net847),
    .X(net306));
 sky130_fd_sc_hd__mux4_1 c374 (.A0(net57),
    .A1(clknet_1_1__leaf_net196),
    .A2(clknet_1_0__leaf_net871),
    .A3(clknet_1_1__leaf_net831),
    .S0(net841),
    .S1(net661),
    .X(net307));
 sky130_fd_sc_hd__mux4_1 c375 (.A0(net193),
    .A1(net167),
    .A2(clknet_1_0__leaf_net871),
    .A3(net905),
    .S0(clknet_1_0__leaf_net196),
    .S1(net847),
    .X(net308));
 sky130_fd_sc_hd__mux4_1 c376 (.A0(net186),
    .A1(net164),
    .A2(net841),
    .A3(clknet_1_0__leaf_net871),
    .S0(net853),
    .S1(net673),
    .X(net309));
 sky130_fd_sc_hd__mux4_1 c377 (.A0(net807),
    .A1(net779),
    .A2(clknet_1_0__leaf_net831),
    .A3(net833),
    .S0(net828),
    .S1(net674),
    .X(net861));
 sky130_fd_sc_hd__xnor2_4 c378 (.A(net80),
    .B(net210),
    .Y(net310));
 sky130_fd_sc_hd__a41o_4 c379 (.A1(net906),
    .A2(net883),
    .A3(net765),
    .A4(net198),
    .B1(net662),
    .X(net311));
 sky130_fd_sc_hd__xnor2_1 c380 (.A(net75),
    .B(net310),
    .Y(net312));
 sky130_fd_sc_hd__xnor2_4 c381 (.A(net201),
    .B(net896),
    .Y(net313));
 sky130_fd_sc_hd__xnor2_2 c382 (.A(net761),
    .B(net82),
    .Y(net314));
 sky130_fd_sc_hd__dfbbp_1 c383 (.CLK(clknet_leaf_40_clk),
    .D(net312),
    .RESET_B(net313),
    .SET_B(net894),
    .Q(net316),
    .Q_N(net315));
 sky130_fd_sc_hd__dfrtp_4 c384 (.CLK(clknet_leaf_40_clk),
    .D(net210),
    .RESET_B(net312),
    .Q(net317));
 sky130_fd_sc_hd__xnor2_4 c385 (.A(net765),
    .B(net317),
    .Y(net318));
 sky130_fd_sc_hd__xnor2_4 c386 (.A(net883),
    .B(net318),
    .Y(net319));
 sky130_fd_sc_hd__xnor2_4 c387 (.A(net894),
    .B(net215),
    .Y(net320));
 sky130_fd_sc_hd__sdfxbp_1 c388 (.CLK(clknet_leaf_40_clk),
    .D(net1000),
    .SCD(net319),
    .SCE(net311),
    .Q(net322),
    .Q_N(net321));
 sky130_fd_sc_hd__xnor2_2 c389 (.A(net313),
    .B(net317),
    .Y(net323));
 sky130_fd_sc_hd__sdfrtp_1 c390 (.CLK(clknet_leaf_40_clk),
    .D(net974),
    .RESET_B(net956),
    .SCD(net319),
    .SCE(net894),
    .Q(net324));
 sky130_fd_sc_hd__dfsbp_1 c391 (.CLK(clknet_leaf_40_clk),
    .D(net951),
    .SET_B(net312),
    .Q(net326),
    .Q_N(net325));
 sky130_fd_sc_hd__sdfxbp_1 c392 (.CLK(clknet_leaf_40_clk),
    .D(net1000),
    .SCD(net311),
    .SCE(net894),
    .Q(net328),
    .Q_N(net327));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net326),
    .A1(net320),
    .A2(net311),
    .A3(net319),
    .S0(net313),
    .S1(net894),
    .X(net329));
 sky130_fd_sc_hd__xnor2_1 c394 (.A(net323),
    .B(net327),
    .Y(net330));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net318),
    .A1(net320),
    .A2(net210),
    .A3(net319),
    .S0(net324),
    .S1(net675),
    .X(net331));
 sky130_fd_sc_hd__sdfxtp_1 c396 (.CLK(clknet_leaf_40_clk),
    .D(net311),
    .SCD(net971),
    .SCE(net676),
    .Q(net332));
 sky130_fd_sc_hd__mux4_1 c397 (.A0(net324),
    .A1(net330),
    .A2(net315),
    .A3(net883),
    .S0(net317),
    .S1(net676),
    .X(net333));
 sky130_fd_sc_hd__mux4_1 c398 (.A0(net328),
    .A1(net332),
    .A2(net333),
    .A3(net883),
    .S0(net916),
    .S1(net676),
    .X(net334));
 sky130_fd_sc_hd__xnor2_1 c399 (.A(net816),
    .B(net310),
    .Y(net335));
 sky130_fd_sc_hd__dfsbp_1 c400 (.CLK(clknet_leaf_37_clk),
    .D(net217),
    .SET_B(net313),
    .Q(net337),
    .Q_N(net336));
 sky130_fd_sc_hd__xnor2_1 c401 (.A(net230),
    .B(net313),
    .Y(net338));
 sky130_fd_sc_hd__sdfrtp_4 c402 (.CLK(clknet_leaf_41_clk),
    .D(net335),
    .RESET_B(net896),
    .SCD(net227),
    .SCE(net229),
    .Q(net339));
 sky130_fd_sc_hd__sdfxtp_2 c403 (.CLK(clknet_leaf_33_clk),
    .D(net333),
    .SCD(net230),
    .SCE(net795),
    .Q(net340));
 sky130_fd_sc_hd__mux4_1 c404 (.A0(net780),
    .A1(net919),
    .A2(net231),
    .A3(net69),
    .S0(net215),
    .S1(net313),
    .X(net341));
 sky130_fd_sc_hd__a21bo_1 c405 (.A1(net340),
    .A2(net816),
    .B1_N(net678),
    .X(net342));
 sky130_fd_sc_hd__mux4_1 c406 (.A0(net335),
    .A1(net232),
    .A2(net340),
    .A3(net101),
    .S0(net336),
    .S1(net678),
    .X(net343));
 sky130_fd_sc_hd__sdfsbp_1 c407 (.CLK(clknet_leaf_38_clk),
    .D(net230),
    .SCD(net340),
    .SCE(net228),
    .SET_B(net943),
    .Q(net345),
    .Q_N(net344));
 sky130_fd_sc_hd__sdfxtp_1 c408 (.CLK(clknet_leaf_38_clk),
    .D(net967),
    .SCD(net335),
    .SCE(net959),
    .Q(net346));
 sky130_fd_sc_hd__xnor2_2 c409 (.A(net346),
    .B(net337),
    .Y(net347));
 sky130_fd_sc_hd__a21bo_2 c410 (.A1(net95),
    .A2(net347),
    .B1_N(net907),
    .X(net348));
 sky130_fd_sc_hd__dfstp_1 c411 (.CLK(clknet_leaf_37_clk),
    .D(net231),
    .SET_B(net944),
    .Q(net349));
 sky130_fd_sc_hd__dfstp_1 c412 (.CLK(clknet_leaf_37_clk),
    .D(net957),
    .SET_B(net319),
    .Q(net350));
 sky130_fd_sc_hd__a21bo_1 c413 (.A1(net101),
    .A2(net84),
    .B1_N(net349),
    .X(net351));
 sky130_fd_sc_hd__a31o_1 c414 (.A1(net337),
    .A2(net101),
    .A3(net350),
    .B1(net313),
    .X(net352));
 sky130_fd_sc_hd__mux4_1 c415 (.A0(net352),
    .A1(net339),
    .A2(net348),
    .A3(net340),
    .S0(net347),
    .S1(net894),
    .X(net353));
 sky130_fd_sc_hd__a21bo_1 c416 (.A1(net353),
    .A2(net350),
    .B1_N(net352),
    .X(net354));
 sky130_fd_sc_hd__a31o_2 c417 (.A1(net345),
    .A2(net354),
    .A3(net350),
    .B1(net347),
    .X(net355));
 sky130_fd_sc_hd__xnor2_4 c418 (.A(net340),
    .B(net677),
    .Y(net356));
 sky130_fd_sc_hd__mux4_1 c419 (.A0(net198),
    .A1(net352),
    .A2(net311),
    .A3(net356),
    .S0(net350),
    .S1(net677),
    .X(net357));
 sky130_fd_sc_hd__xnor2_4 c420 (.A(net98),
    .B(net680),
    .Y(net358));
 sky130_fd_sc_hd__a21bo_1 c421 (.A1(net100),
    .A2(net215),
    .B1_N(net885),
    .X(net359));
 sky130_fd_sc_hd__a21bo_1 c422 (.A1(net354),
    .A2(net359),
    .B1_N(net896),
    .X(net842));
 sky130_fd_sc_hd__sdfsbp_1 c423 (.CLK(clknet_leaf_2_clk),
    .D(net347),
    .SCD(net880),
    .SCE(net224),
    .SET_B(net354),
    .Q(net361),
    .Q_N(net360));
 sky130_fd_sc_hd__mux4_1 c424 (.A0(net351),
    .A1(net265),
    .A2(net311),
    .A3(net251),
    .S0(net880),
    .S1(clknet_1_0__leaf_net859),
    .X(net362));
 sky130_fd_sc_hd__dfbbn_1 c425 (.CLK_N(clknet_leaf_37_clk),
    .D(net224),
    .RESET_B(net228),
    .SET_B(net682),
    .Q(net364),
    .Q_N(net363));
 sky130_fd_sc_hd__sdfbbn_1 c426 (.CLK_N(clknet_leaf_37_clk),
    .D(net811),
    .RESET_B(net963),
    .SCD(net234),
    .SCE(net311),
    .SET_B(net900),
    .Q(net839),
    .Q_N(net365));
 sky130_fd_sc_hd__a21bo_1 c427 (.A1(net358),
    .A2(net224),
    .B1_N(net365),
    .X(net366));
 sky130_fd_sc_hd__dfbbn_2 c428 (.CLK_N(clknet_leaf_2_clk),
    .D(net0),
    .RESET_B(net100),
    .SET_B(net311),
    .Q(net368),
    .Q_N(net367));
 sky130_fd_sc_hd__sdfstp_1 c429 (.CLK(clknet_leaf_2_clk),
    .D(net310),
    .SCD(net251),
    .SCE(net802),
    .SET_B(net367),
    .Q(net369));
 sky130_fd_sc_hd__a31o_2 c430 (.A1(net364),
    .A2(net234),
    .A3(net367),
    .B1(net369),
    .X(net370));
 sky130_fd_sc_hd__a41o_1 c431 (.A1(net350),
    .A2(net366),
    .A3(net105),
    .A4(net355),
    .B1(net370),
    .X(net371));
 sky130_fd_sc_hd__a41o_4 c432 (.A1(net366),
    .A2(net370),
    .A3(net368),
    .A4(net358),
    .B1(net811),
    .X(net372));
 sky130_fd_sc_hd__a31o_2 c433 (.A1(net369),
    .A2(net347),
    .A3(net367),
    .B1(net372),
    .X(net844));
 sky130_fd_sc_hd__a41o_1 c434 (.A1(net105),
    .A2(net839),
    .A3(net761),
    .A4(net310),
    .B1(clknet_1_1__leaf_net130),
    .X(net373));
 sky130_fd_sc_hd__mux4_1 c435 (.A0(net340),
    .A1(net350),
    .A2(net358),
    .A3(net310),
    .S0(net844),
    .S1(net370),
    .X(net374));
 sky130_fd_sc_hd__a41o_1 c436 (.A1(net372),
    .A2(net358),
    .A3(net367),
    .A4(clknet_1_0__leaf_net130),
    .B1(net683),
    .X(net375));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(net359),
    .A1(clknet_1_0__leaf_net375),
    .A2(net98),
    .A3(net105),
    .S0(net681),
    .S1(net683),
    .X(net376));
 sky130_fd_sc_hd__sdfstp_2 c438 (.CLK(clknet_leaf_35_clk),
    .D(net368),
    .SCD(clknet_1_1__leaf_net373),
    .SCE(net908),
    .SET_B(net249),
    .Q(net377));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net377),
    .A1(net368),
    .A2(clknet_1_0__leaf_net373),
    .A3(net372),
    .S0(net370),
    .S1(net1002),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 c440 (.A0(net844),
    .A1(net377),
    .A2(net310),
    .A3(net679),
    .S0(net1002),
    .S1(net999),
    .X(net379));
 sky130_fd_sc_hd__dfbbp_1 c441 (.CLK(clknet_leaf_4_clk),
    .D(net249),
    .RESET_B(net358),
    .SET_B(net265),
    .Q(net381),
    .Q_N(net380));
 sky130_fd_sc_hd__a21bo_1 c442 (.A1(net792),
    .A2(net380),
    .B1_N(net668),
    .X(net382));
 sky130_fd_sc_hd__a21bo_1 c443 (.A1(net785),
    .A2(net265),
    .B1_N(clknet_1_0__leaf_net655),
    .X(net383));
 sky130_fd_sc_hd__a21bo_2 c444 (.A1(net802),
    .A2(net151),
    .B1_N(net761),
    .X(net851));
 sky130_fd_sc_hd__mux4_1 c445 (.A0(net884),
    .A1(net770),
    .A2(net851),
    .A3(net844),
    .S0(net21),
    .S1(net665),
    .X(net384));
 sky130_fd_sc_hd__sdfxbp_1 c446 (.CLK(clknet_leaf_24_clk),
    .D(net908),
    .SCD(clknet_1_1__leaf_net281),
    .SCE(clknet_1_1__leaf_net686),
    .Q(net873),
    .Q_N(net385));
 sky130_fd_sc_hd__a21bo_1 c447 (.A1(net894),
    .A2(net274),
    .B1_N(clknet_1_1__leaf_net654),
    .X(net855));
 sky130_fd_sc_hd__a31o_1 c448 (.A1(net887),
    .A2(net21),
    .A3(net904),
    .B1(clknet_1_0__leaf_net687),
    .X(net386));
 sky130_fd_sc_hd__sdfxbp_1 c449 (.CLK(clknet_leaf_14_clk),
    .D(net381),
    .SCD(clknet_1_0__leaf_net281),
    .SCE(clknet_1_0__leaf_net386),
    .Q(net388),
    .Q_N(net387));
 sky130_fd_sc_hd__a31o_1 c450 (.A1(net370),
    .A2(net388),
    .A3(net907),
    .B1(clknet_1_0__leaf_net386),
    .X(net389));
 sky130_fd_sc_hd__sdfbbp_1 c451 (.CLK(clknet_leaf_3_clk),
    .D(net266),
    .RESET_B(clknet_1_0__leaf_net386),
    .SCD(net274),
    .SCE(net987),
    .SET_B(net802),
    .Q(net391),
    .Q_N(net390));
 sky130_fd_sc_hd__mux4_1 c452 (.A0(net265),
    .A1(net371),
    .A2(clknet_1_0__leaf_net386),
    .A3(net356),
    .S0(clknet_1_1__leaf_net389),
    .S1(net377),
    .X(net392));
 sky130_fd_sc_hd__a41o_1 c453 (.A1(net215),
    .A2(net390),
    .A3(clknet_1_0__leaf_net386),
    .A4(net904),
    .B1(net665),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 c454 (.A0(net383),
    .A1(net372),
    .A2(clknet_1_0__leaf_net855),
    .A3(net832),
    .S0(clknet_1_0__leaf_net393),
    .S1(net390),
    .X(net394));
 sky130_fd_sc_hd__a41o_1 c455 (.A1(net387),
    .A2(clknet_1_1__leaf_net389),
    .A3(clknet_1_0__leaf_net386),
    .A4(net274),
    .B1(net688),
    .X(net826));
 sky130_fd_sc_hd__sdfxtp_1 c456 (.CLK(clknet_leaf_11_clk),
    .D(net382),
    .SCD(clknet_1_1__leaf_net826),
    .SCE(clknet_1_1__leaf_net859),
    .Q(net849));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(net361),
    .A1(net851),
    .A2(clknet_1_1__leaf_net389),
    .A3(net387),
    .S0(net668),
    .S1(net689),
    .X(net395));
 sky130_fd_sc_hd__a21bo_1 c458 (.A1(clknet_1_1__leaf_net154),
    .A2(clknet_1_0__leaf_net686),
    .B1_N(clknet_1_0__leaf_net687),
    .X(net396));
 sky130_fd_sc_hd__a21bo_1 c459 (.A1(clknet_1_1__leaf_net393),
    .A2(net274),
    .B1_N(clknet_1_0__leaf_net386),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net397),
    .A1(net13),
    .A2(net360),
    .A3(net370),
    .S0(net265),
    .S1(net887),
    .X(net398));
 sky130_fd_sc_hd__a41o_1 c461 (.A1(net396),
    .A2(clknet_1_0__leaf_net855),
    .A3(clknet_1_0__leaf_net386),
    .A4(net904),
    .B1(net900),
    .X(net399));
 sky130_fd_sc_hd__sdfbbn_1 c462 (.CLK_N(clknet_leaf_13_clk),
    .D(net300),
    .RESET_B(net887),
    .SCD(net288),
    .SCE(net28),
    .SET_B(clknet_1_0__leaf_net671),
    .Q(net401),
    .Q_N(net400));
 sky130_fd_sc_hd__mux4_1 c463 (.A0(net395),
    .A1(net300),
    .A2(net897),
    .A3(net296),
    .S0(net28),
    .S1(clknet_1_1__leaf_net655),
    .X(net402));
 sky130_fd_sc_hd__mux4_1 c464 (.A0(net293),
    .A1(net289),
    .A2(net851),
    .A3(net28),
    .S0(clknet_1_0__leaf_net671),
    .S1(clknet_1_0__leaf_net672),
    .X(net403));
 sky130_fd_sc_hd__a41o_1 c465 (.A1(net297),
    .A2(clknet_1_1__leaf_net855),
    .A3(net884),
    .A4(net289),
    .B1(net875),
    .X(net404));
 sky130_fd_sc_hd__a41o_1 c466 (.A1(net291),
    .A2(net28),
    .A3(clknet_1_0__leaf_net386),
    .A4(net679),
    .B1(clknet_1_1__leaf_net687),
    .X(net846));
 sky130_fd_sc_hd__sdfbbn_1 c467 (.CLK_N(clknet_leaf_15_clk),
    .D(net169),
    .RESET_B(net897),
    .SCD(net908),
    .SCE(clknet_1_1__leaf_net404),
    .SET_B(net12),
    .Q(net405));
 sky130_fd_sc_hd__mux4_1 c468 (.A0(net28),
    .A1(net852),
    .A2(net832),
    .A3(net884),
    .S0(clknet_1_0__leaf_net404),
    .S1(net905),
    .X(net406));
 sky130_fd_sc_hd__a41o_1 c469 (.A1(net885),
    .A2(net28),
    .A3(net851),
    .A4(clknet_1_0__leaf_net386),
    .B1(net694),
    .X(net407));
 sky130_fd_sc_hd__sdfbbp_1 c470 (.CLK(clknet_leaf_14_clk),
    .D(net401),
    .RESET_B(net368),
    .SCD(clknet_1_0__leaf_net404),
    .SCE(net289),
    .SET_B(net953),
    .Q(net409),
    .Q_N(net408));
 sky130_fd_sc_hd__mux4_1 c471 (.A0(net289),
    .A1(clknet_1_0__leaf_net846),
    .A2(net300),
    .A3(net887),
    .S0(clknet_1_1__leaf_net671),
    .S1(clknet_1_1__leaf_net687),
    .X(net410));
 sky130_fd_sc_hd__sdfbbn_1 c472 (.CLK_N(clknet_leaf_14_clk),
    .D(clknet_1_0__leaf_net404),
    .RESET_B(net964),
    .SCD(net409),
    .SCE(net224),
    .SET_B(net975),
    .Q(net843));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(net388),
    .A1(net300),
    .A2(net408),
    .A3(net291),
    .S0(clknet_1_1__leaf_net859),
    .S1(net848),
    .X(net411));
 sky130_fd_sc_hd__sdfbbn_1 c474 (.CLK_N(clknet_leaf_12_clk),
    .D(net358),
    .RESET_B(clknet_1_1__leaf_net404),
    .SCD(net888),
    .SCE(net905),
    .SET_B(net860),
    .Q(net413),
    .Q_N(net412));
 sky130_fd_sc_hd__a41o_1 c475 (.A1(net287),
    .A2(net388),
    .A3(clknet_1_0__leaf_net386),
    .A4(clknet_1_1__leaf_net859),
    .B1(net860),
    .X(net856));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(net413),
    .A1(net289),
    .A2(net904),
    .A3(net850),
    .S0(clknet_1_0__leaf_net826),
    .S1(net365),
    .X(net414));
 sky130_fd_sc_hd__a41o_1 c477 (.A1(net850),
    .A2(clknet_1_0__leaf_net403),
    .A3(net412),
    .A4(net693),
    .B1(net695),
    .X(net415));
 sky130_fd_sc_hd__a41o_1 c478 (.A1(net409),
    .A2(net413),
    .A3(clknet_1_0__leaf_net386),
    .A4(net904),
    .B1(net694),
    .X(net416));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(net288),
    .A1(net413),
    .A2(net291),
    .A3(clknet_1_1__leaf_net859),
    .S0(net679),
    .S1(net695),
    .X(net417));
 sky130_fd_sc_hd__sdfbbp_1 c480 (.CLK(clknet_leaf_18_clk),
    .D(net405),
    .RESET_B(net417),
    .SCD(net905),
    .SCE(clknet_1_0__leaf_net826),
    .SET_B(net694),
    .Q(net840));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net407),
    .A1(net416),
    .A2(net851),
    .A3(net169),
    .S0(net412),
    .S1(net694),
    .X(net418));
 sky130_fd_sc_hd__sdfbbn_1 c482 (.CLK_N(clknet_leaf_17_clk),
    .D(net887),
    .RESET_B(net415),
    .SCD(net412),
    .SCE(net692),
    .SET_B(net858),
    .Q(net420),
    .Q_N(net419));
 sky130_fd_sc_hd__xnor2_4 c504 (.A(net82),
    .B(net675),
    .Y(net421));
 sky130_fd_sc_hd__xnor2_1 c505 (.A(net819),
    .B(net84),
    .Y(net422));
 sky130_fd_sc_hd__xnor2_4 c506 (.A(net891),
    .B(net421),
    .Y(net423));
 sky130_fd_sc_hd__xnor2_4 c507 (.A(net936),
    .B(net332),
    .Y(net424));
 sky130_fd_sc_hd__xnor2_4 c508 (.A(net916),
    .B(net320),
    .Y(net425));
 sky130_fd_sc_hd__xnor2_1 c509 (.A(net216),
    .B(net924),
    .Y(net426));
 sky130_fd_sc_hd__a21bo_4 c510 (.A1(net425),
    .A2(net891),
    .B1_N(net916),
    .X(net427));
 sky130_fd_sc_hd__sdfxtp_1 c511 (.CLK(clknet_leaf_32_clk),
    .D(net323),
    .SCD(net333),
    .SCE(net889),
    .Q(net428));
 sky130_fd_sc_hd__sdfxtp_4 c512 (.CLK(clknet_leaf_32_clk),
    .D(net889),
    .SCD(net319),
    .SCE(net425),
    .Q(net837));
 sky130_fd_sc_hd__dfbbn_1 c513 (.CLK_N(clknet_leaf_33_clk),
    .D(net426),
    .RESET_B(net891),
    .SET_B(net427),
    .Q(net430),
    .Q_N(net429));
 sky130_fd_sc_hd__xnor2_4 c514 (.A(net425),
    .B(net889),
    .Y(net431));
 sky130_fd_sc_hd__xnor2_4 c515 (.A(net937),
    .B(net837),
    .Y(net432));
 sky130_fd_sc_hd__a21bo_1 c516 (.A1(net431),
    .A2(net890),
    .B1_N(net891),
    .X(net433));
 sky130_fd_sc_hd__dfbbn_1 c517 (.CLK_N(clknet_leaf_32_clk),
    .D(net977),
    .RESET_B(net426),
    .SET_B(net318),
    .Q(net435),
    .Q_N(net434));
 sky130_fd_sc_hd__xnor2_4 c518 (.A(net424),
    .B(net206),
    .Y(net436));
 sky130_fd_sc_hd__mux4_1 c519 (.A0(net435),
    .A1(net427),
    .A2(net436),
    .A3(net425),
    .S0(net431),
    .S1(net432),
    .X(net437));
 sky130_fd_sc_hd__mux4_2 c520 (.A0(net434),
    .A1(net317),
    .A2(net436),
    .A3(net837),
    .S0(net427),
    .S1(net891),
    .X(net438));
 sky130_fd_sc_hd__a41o_1 c521 (.A1(net928),
    .A2(net431),
    .A3(net772),
    .A4(net892),
    .B1(net662),
    .X(net439));
 sky130_fd_sc_hd__mux4_2 c522 (.A0(net433),
    .A1(net437),
    .A2(net428),
    .A3(net427),
    .S0(net895),
    .S1(net891),
    .X(net440));
 sky130_fd_sc_hd__mux4_1 c523 (.A0(net427),
    .A1(net425),
    .A2(net881),
    .A3(net925),
    .S0(net931),
    .S1(net894),
    .X(net441));
 sky130_fd_sc_hd__dfbbp_1 c524 (.CLK(clknet_leaf_31_clk),
    .D(net441),
    .RESET_B(net926),
    .SET_B(net71),
    .Q(net442));
 sky130_fd_sc_hd__a21bo_1 c525 (.A1(net342),
    .A2(net431),
    .B1_N(net891),
    .X(net443));
 sky130_fd_sc_hd__xnor2_4 c526 (.A(net919),
    .B(net832),
    .Y(net444));
 sky130_fd_sc_hd__xnor2_1 c527 (.A(net431),
    .B(net355),
    .Y(net445));
 sky130_fd_sc_hd__a21bo_1 c528 (.A1(net84),
    .A2(net885),
    .B1_N(net423),
    .X(net446));
 sky130_fd_sc_hd__dfstp_2 c529 (.CLK(clknet_leaf_33_clk),
    .D(net426),
    .SET_B(net446),
    .Q(net447));
 sky130_fd_sc_hd__xnor2_1 c530 (.A(net330),
    .B(net432),
    .Y(net448));
 sky130_fd_sc_hd__a21bo_1 c531 (.A1(net447),
    .A2(net84),
    .B1_N(net355),
    .X(net449));
 sky130_fd_sc_hd__a21bo_4 c532 (.A1(net438),
    .A2(net978),
    .B1_N(net891),
    .X(net450));
 sky130_fd_sc_hd__mux4_1 c533 (.A0(net449),
    .A1(net233),
    .A2(net447),
    .A3(net348),
    .S0(net227),
    .S1(net879),
    .X(net451));
 sky130_fd_sc_hd__a21bo_4 c534 (.A1(net338),
    .A2(net69),
    .B1_N(net423),
    .X(net452));
 sky130_fd_sc_hd__xnor2_1 c535 (.A(net892),
    .B(net339),
    .Y(net453));
 sky130_fd_sc_hd__xnor2_1 c536 (.A(net450),
    .B(net313),
    .Y(net454));
 sky130_fd_sc_hd__a41o_2 c537 (.A1(net227),
    .A2(net825),
    .A3(net793),
    .A4(net881),
    .B1(net985),
    .X(net455));
 sky130_fd_sc_hd__mux4_1 c538 (.A0(net445),
    .A1(net452),
    .A2(net932),
    .A3(net879),
    .S0(net348),
    .S1(net770),
    .X(net456));
 sky130_fd_sc_hd__sdfstp_1 c539 (.CLK(clknet_leaf_33_clk),
    .D(net319),
    .SCD(net448),
    .SCE(net452),
    .SET_B(net450),
    .Q(net457));
 sky130_fd_sc_hd__sdfbbn_1 c540 (.CLK_N(clknet_2_0__leaf_clk),
    .D(net448),
    .RESET_B(net447),
    .SCD(net455),
    .SCE(net445),
    .SET_B(net319),
    .Q(net459),
    .Q_N(net458));
 sky130_fd_sc_hd__mux4_1 c541 (.A0(net453),
    .A1(net450),
    .A2(net927),
    .A3(net452),
    .S0(net444),
    .S1(net459),
    .X(net460));
 sky130_fd_sc_hd__mux4_1 c542 (.A0(net457),
    .A1(net779),
    .A2(net338),
    .A3(net313),
    .S0(net447),
    .S1(net348),
    .X(net461));
 sky130_fd_sc_hd__sdfbbp_1 c543 (.CLK(clknet_leaf_33_clk),
    .D(net461),
    .RESET_B(net455),
    .SCD(net432),
    .SCE(net431),
    .SET_B(net947),
    .Q(net463),
    .Q_N(net462));
 sky130_fd_sc_hd__sdfbbn_2 c544 (.CLK_N(clknet_leaf_33_clk),
    .D(net446),
    .RESET_B(net892),
    .SCD(net461),
    .SCE(net449),
    .SET_B(net699),
    .Q(net465),
    .Q_N(net464));
 sky130_fd_sc_hd__mux4_1 c545 (.A0(net214),
    .A1(net935),
    .A2(net453),
    .A3(net465),
    .S0(net792),
    .S1(net458),
    .X(net466));
 sky130_fd_sc_hd__dlrbn_1 c546 (.D(net896),
    .GATE_N(clknet_leaf_35_clk),
    .RESET_B(net879),
    .Q(net468),
    .Q_N(net467));
 sky130_fd_sc_hd__dlrbn_1 c547 (.D(net311),
    .GATE_N(clknet_leaf_35_clk),
    .RESET_B(net978),
    .Q(net470),
    .Q_N(net469));
 sky130_fd_sc_hd__xnor2_1 c548 (.A(net469),
    .B(net958),
    .Y(net471));
 sky130_fd_sc_hd__a21bo_2 c549 (.A1(net355),
    .A2(net459),
    .B1_N(net934),
    .X(net472));
 sky130_fd_sc_hd__dlrbp_1 c550 (.D(clknet_1_1__leaf_net375),
    .GATE(clknet_leaf_35_clk),
    .RESET_B(net950),
    .Q(net473));
 sky130_fd_sc_hd__xnor2_4 c551 (.A(net800),
    .B(net355),
    .Y(net474));
 sky130_fd_sc_hd__a21bo_2 c552 (.A1(net471),
    .A2(net450),
    .B1_N(net981),
    .X(net475));
 sky130_fd_sc_hd__a21bo_2 c553 (.A1(net459),
    .A2(net470),
    .B1_N(net800),
    .X(net476));
 sky130_fd_sc_hd__dlrbp_1 c554 (.D(net474),
    .GATE(clknet_leaf_25_clk),
    .RESET_B(net1004),
    .Q(net477));
 sky130_fd_sc_hd__a21bo_1 c555 (.A1(net795),
    .A2(net476),
    .B1_N(net452),
    .X(net478));
 sky130_fd_sc_hd__sdfxbp_1 c556 (.CLK(clknet_leaf_36_clk),
    .D(clknet_1_1__leaf_net130),
    .SCD(net472),
    .SCE(net262),
    .Q(net479));
 sky130_fd_sc_hd__dlrtn_1 c557 (.D(net454),
    .GATE_N(clknet_leaf_34_clk),
    .RESET_B(net947),
    .Q(net480));
 sky130_fd_sc_hd__a21bo_2 c558 (.A1(net477),
    .A2(net480),
    .B1_N(net377),
    .X(net829));
 sky130_fd_sc_hd__mux4_1 c559 (.A0(net98),
    .A1(net263),
    .A2(net480),
    .A3(net825),
    .S0(net311),
    .S1(net472),
    .X(net481));
 sky130_fd_sc_hd__a21bo_4 c560 (.A1(net478),
    .A2(net480),
    .B1_N(net701),
    .X(net482));
 sky130_fd_sc_hd__xnor2_1 c561 (.A(net482),
    .B(net701),
    .Y(net483));
 sky130_fd_sc_hd__a31o_1 c562 (.A1(net473),
    .A2(net467),
    .A3(net881),
    .B1(net701),
    .X(net484));
 sky130_fd_sc_hd__a31o_1 c563 (.A1(net470),
    .A2(net476),
    .A3(net837),
    .B1(net701),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c564 (.A0(net480),
    .A1(net997),
    .A2(net482),
    .A3(net880),
    .S0(net484),
    .S1(net485),
    .X(net486));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net483),
    .A1(net450),
    .A2(net485),
    .A3(net98),
    .S0(net908),
    .S1(clknet_1_0__leaf_net702),
    .X(net487));
 sky130_fd_sc_hd__sdfbbn_1 c566 (.CLK_N(clknet_leaf_34_clk),
    .D(net263),
    .RESET_B(net487),
    .SCD(net443),
    .SCE(net476),
    .SET_B(clknet_1_1__leaf_net702),
    .Q(net488));
 sky130_fd_sc_hd__a31o_1 c567 (.A1(net391),
    .A2(net377),
    .A3(net465),
    .B1(net980),
    .X(net489));
 sky130_fd_sc_hd__sedfxbp_1 c568 (.CLK(clknet_leaf_15_clk),
    .D(net484),
    .DE(net881),
    .SCD(net485),
    .SCE(clknet_1_0__leaf_net281),
    .Q(net490));
 sky130_fd_sc_hd__a41o_1 c569 (.A1(net894),
    .A2(net485),
    .A3(net884),
    .A4(net150),
    .B1(net669),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net356),
    .A1(net472),
    .A2(net908),
    .A3(net391),
    .S0(net228),
    .S1(clknet_1_0__leaf_net281),
    .X(net492));
 sky130_fd_sc_hd__sdfbbp_1 c571 (.CLK(clknet_leaf_35_clk),
    .D(net489),
    .RESET_B(net356),
    .SCD(net901),
    .SCE(net467),
    .SET_B(net878),
    .Q(net494),
    .Q_N(net493));
 sky130_fd_sc_hd__sdfbbn_1 c572 (.CLK_N(clknet_leaf_35_clk),
    .D(net452),
    .RESET_B(net217),
    .SCD(clknet_1_0__leaf_net389),
    .SCE(net878),
    .SET_B(clknet_1_1__leaf_net655),
    .Q(net495));
 sky130_fd_sc_hd__a41o_1 c573 (.A1(net468),
    .A2(net452),
    .A3(net894),
    .A4(net897),
    .B1(net356),
    .X(net496));
 sky130_fd_sc_hd__sdfbbn_1 c574 (.CLK_N(clknet_leaf_15_clk),
    .D(net485),
    .RESET_B(net12),
    .SCD(clknet_1_0__leaf_net281),
    .SCE(net377),
    .SET_B(net900),
    .Q(net498),
    .Q_N(net497));
 sky130_fd_sc_hd__mux4_1 c575 (.A0(net228),
    .A1(net825),
    .A2(net476),
    .A3(clknet_1_0__leaf_net389),
    .S0(net497),
    .S1(clknet_1_1__leaf_net386),
    .X(net499));
 sky130_fd_sc_hd__a31o_2 c576 (.A1(net151),
    .A2(net356),
    .A3(net829),
    .B1(net465),
    .X(net500));
 sky130_fd_sc_hd__a31o_1 c577 (.A1(net399),
    .A2(net488),
    .A3(net468),
    .B1(net496),
    .X(net501));
 sky130_fd_sc_hd__sdfbbp_1 c578 (.CLK(clknet_leaf_24_clk),
    .D(net446),
    .RESET_B(net385),
    .SCD(clknet_1_0__leaf_net501),
    .SCE(net906),
    .SET_B(net703),
    .Q(net503),
    .Q_N(net502));
 sky130_fd_sc_hd__mux4_1 c579 (.A0(net476),
    .A1(net496),
    .A2(net493),
    .A3(net502),
    .S0(clknet_1_0__leaf_net501),
    .S1(net900),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c580 (.A0(clknet_1_0__leaf_net389),
    .A1(net446),
    .A2(net468),
    .A3(net503),
    .S0(net476),
    .S1(clknet_1_1__leaf_net655),
    .X(net505));
 sky130_fd_sc_hd__sdfbbn_1 c581 (.CLK_N(clknet_leaf_23_clk),
    .D(net969),
    .RESET_B(net377),
    .SCD(net837),
    .SCE(clknet_1_1__leaf_net501),
    .SET_B(net502),
    .Q(net506));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(net506),
    .A1(net500),
    .A2(net377),
    .A3(clknet_1_1__leaf_net501),
    .S0(net502),
    .S1(clknet_1_0__leaf_net834),
    .X(net507));
 sky130_fd_sc_hd__sdfbbn_1 c583 (.CLK_N(clknet_leaf_24_clk),
    .D(net968),
    .RESET_B(net494),
    .SCD(net500),
    .SCE(net503),
    .SET_B(net475),
    .Q(net509),
    .Q_N(net508));
 sky130_fd_sc_hd__mux4_1 c584 (.A0(clknet_1_0__leaf_net501),
    .A1(net505),
    .A2(net508),
    .A3(net895),
    .S0(net912),
    .S1(net476),
    .X(net510));
 sky130_fd_sc_hd__a31o_1 c585 (.A1(net503),
    .A2(net476),
    .A3(net704),
    .B1(net705),
    .X(net511));
 sky130_fd_sc_hd__sdfbbp_1 c586 (.CLK(clknet_leaf_23_clk),
    .D(net371),
    .RESET_B(net511),
    .SCD(net825),
    .SCE(net502),
    .SET_B(clknet_1_1__leaf_net501),
    .Q(net512));
 sky130_fd_sc_hd__sdfbbn_1 c587 (.CLK_N(clknet_leaf_23_clk),
    .D(net970),
    .RESET_B(net503),
    .SCD(clknet_1_1__leaf_net501),
    .SCE(net511),
    .SET_B(net837),
    .Q(net513));
 sky130_fd_sc_hd__sdfbbn_1 c588 (.CLK_N(clknet_leaf_23_clk),
    .D(net224),
    .RESET_B(net888),
    .SCD(net462),
    .SCE(clknet_1_0__leaf_net826),
    .SET_B(net822),
    .Q(net515),
    .Q_N(net514));
 sky130_fd_sc_hd__sdfbbp_1 c589 (.CLK(clknet_leaf_15_clk),
    .D(net420),
    .RESET_B(net772),
    .SCD(net913),
    .SCE(net224),
    .SET_B(net829),
    .Q(net517),
    .Q_N(net516));
 sky130_fd_sc_hd__sdfbbn_1 c590 (.CLK_N(clknet_leaf_15_clk),
    .D(net472),
    .RESET_B(net517),
    .SCD(net829),
    .SCE(clknet_1_0__leaf_net299),
    .SET_B(net695),
    .Q(net518));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(net12),
    .A1(clknet_1_0__leaf_net299),
    .A2(net908),
    .A3(clknet_1_0__leaf_net826),
    .S0(net779),
    .S1(net695),
    .X(net519));
 sky130_fd_sc_hd__mux4_1 c592 (.A0(net513),
    .A1(net516),
    .A2(net888),
    .A3(clknet_1_0__leaf_net826),
    .S0(net694),
    .S1(clknet_1_1__leaf_net834),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(clknet_1_1__leaf_net299),
    .A1(net464),
    .A2(net372),
    .A3(net691),
    .S0(net693),
    .S1(net694),
    .X(net521));
 sky130_fd_sc_hd__sdfbbn_1 c594 (.CLK_N(clknet_leaf_22_clk),
    .D(clknet_1_1__leaf_net299),
    .RESET_B(net372),
    .SCD(net514),
    .SCE(net888),
    .SET_B(net960),
    .Q(net523),
    .Q_N(net522));
 sky130_fd_sc_hd__sdfbbp_1 c595 (.CLK(clknet_leaf_16_clk),
    .D(net880),
    .RESET_B(net888),
    .SCD(clknet_1_1__leaf_net655),
    .SCE(net984),
    .SET_B(net708),
    .Q(net525),
    .Q_N(net524));
 sky130_fd_sc_hd__a41o_1 c596 (.A1(net524),
    .A2(net882),
    .A3(net706),
    .A4(net707),
    .B1(net708),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 c597 (.A0(net463),
    .A1(net512),
    .A2(net829),
    .A3(clknet_1_1__leaf_net655),
    .S0(net695),
    .S1(net708),
    .X(net527));
 sky130_fd_sc_hd__mux4_1 c598 (.A0(net490),
    .A1(net420),
    .A2(net837),
    .A3(net464),
    .S0(net900),
    .S1(net695),
    .X(net528));
 sky130_fd_sc_hd__mux4_1 c599 (.A0(net518),
    .A1(net792),
    .A2(net825),
    .A3(net879),
    .S0(clknet_1_1__leaf_net655),
    .S1(net706),
    .X(net529));
 sky130_fd_sc_hd__a41o_1 c600 (.A1(net527),
    .A2(net837),
    .A3(net694),
    .A4(net708),
    .B1(net709),
    .X(net530));
 sky130_fd_sc_hd__mux4_1 c601 (.A0(clknet_1_1__leaf_net403),
    .A1(net528),
    .A2(net837),
    .A3(net875),
    .S0(clknet_1_0__leaf_net834),
    .S1(net708),
    .X(net531));
 sky130_fd_sc_hd__sdfbbn_1 c602 (.CLK_N(clknet_leaf_17_clk),
    .D(clknet_1_0__leaf_net531),
    .RESET_B(net888),
    .SCD(net989),
    .SCE(net298),
    .SET_B(net966),
    .Q(net877),
    .Q_N(net532));
 sky130_fd_sc_hd__mux4_2 c603 (.A0(net884),
    .A1(net532),
    .A2(net875),
    .A3(net706),
    .S0(net707),
    .S1(net709),
    .X(net533));
 sky130_fd_sc_hd__sdfbbn_1 c604 (.CLK_N(clknet_leaf_16_clk),
    .D(net772),
    .RESET_B(net908),
    .SCD(net994),
    .SCE(net533),
    .SET_B(net966),
    .Q(net535),
    .Q_N(net534));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net138),
    .A1(net533),
    .A2(clknet_1_1__leaf_net531),
    .A3(net532),
    .S0(net472),
    .S1(net692),
    .X(net536));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net530),
    .A1(net908),
    .A2(net534),
    .A3(net533),
    .S0(net709),
    .S1(net988),
    .X(net537));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(net525),
    .A1(net877),
    .A2(net535),
    .A3(net779),
    .S0(net533),
    .S1(net988),
    .X(net538));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net534),
    .A1(net690),
    .A2(net695),
    .A3(net708),
    .S0(net710),
    .S1(net712),
    .X(net539));
 sky130_fd_sc_hd__mux4_2 c62 (.A0(net800),
    .A1(net798),
    .A2(net760),
    .A3(net818),
    .S0(net771),
    .S1(net802),
    .X(net0));
 sky130_fd_sc_hd__xnor2_1 c63 (.A(net798),
    .B(net901),
    .Y(net1));
 sky130_fd_sc_hd__xnor2_1 c630 (.A(net71),
    .B(net891),
    .Y(net540));
 sky130_fd_sc_hd__a31o_2 c631 (.A1(net428),
    .A2(net770),
    .A3(net930),
    .B1(net889),
    .X(net541));
 sky130_fd_sc_hd__xnor2_4 c632 (.A(net541),
    .B(net885),
    .Y(net542));
 sky130_fd_sc_hd__xnor2_1 c633 (.A(net541),
    .B(net542),
    .Y(net543));
 sky130_fd_sc_hd__xnor2_4 c634 (.A(net890),
    .B(net917),
    .Y(net544));
 sky130_fd_sc_hd__xnor2_2 c635 (.A(net430),
    .B(net69),
    .Y(net545));
 sky130_fd_sc_hd__dlrtn_1 c636 (.D(net543),
    .GATE_N(clknet_leaf_31_clk),
    .RESET_B(net889),
    .Q(net546));
 sky130_fd_sc_hd__xnor2_1 c637 (.A(net544),
    .B(net542),
    .Y(net547));
 sky130_fd_sc_hd__xnor2_4 c638 (.A(net544),
    .B(net917),
    .Y(net548));
 sky130_fd_sc_hd__a21bo_1 c639 (.A1(net442),
    .A2(net540),
    .B1_N(net891),
    .X(net549));
 sky130_fd_sc_hd__xnor2_4 c64 (.A(net813),
    .B(net4),
    .Y(net2));
 sky130_fd_sc_hd__xnor2_4 c640 (.A(net318),
    .B(net542),
    .Y(net550));
 sky130_fd_sc_hd__xnor2_2 c641 (.A(net548),
    .B(net542),
    .Y(net551));
 sky130_fd_sc_hd__xnor2_1 c642 (.A(net542),
    .B(net918),
    .Y(net552));
 sky130_fd_sc_hd__dlrtn_2 c643 (.D(net546),
    .GATE_N(clknet_leaf_31_clk),
    .RESET_B(net551),
    .Q(net553));
 sky130_fd_sc_hd__mux4_1 c644 (.A0(net549),
    .A1(net546),
    .A2(net553),
    .A3(net551),
    .S0(net548),
    .S1(net892),
    .X(net554));
 sky130_fd_sc_hd__xnor2_2 c645 (.A(net439),
    .B(net553),
    .Y(net555));
 sky130_fd_sc_hd__sedfxbp_1 c646 (.CLK(clknet_leaf_29_clk),
    .D(net551),
    .DE(net881),
    .SCD(net553),
    .SCE(net976),
    .Q(net557),
    .Q_N(net556));
 sky130_fd_sc_hd__a31o_2 c647 (.A1(net553),
    .A2(net556),
    .A3(net892),
    .B1(net713),
    .X(net558));
 sky130_fd_sc_hd__a31o_1 c648 (.A1(net540),
    .A2(net553),
    .A3(net548),
    .B1(net549),
    .X(net559));
 sky130_fd_sc_hd__mux4_1 c649 (.A0(net557),
    .A1(net559),
    .A2(net543),
    .A3(net551),
    .S0(net555),
    .S1(net558),
    .X(net560));
 sky130_fd_sc_hd__xnor2_4 c65 (.A(net820),
    .B(net909),
    .Y(net3));
 sky130_fd_sc_hd__mux4_1 c650 (.A0(net437),
    .A1(net559),
    .A2(net551),
    .A3(net542),
    .S0(net69),
    .S1(net1001),
    .X(net561));
 sky130_fd_sc_hd__a31o_1 c651 (.A1(net232),
    .A2(net317),
    .A3(net339),
    .B1(net464),
    .X(net562));
 sky130_fd_sc_hd__a21bo_1 c652 (.A1(net562),
    .A2(net317),
    .B1_N(net548),
    .X(net563));
 sky130_fd_sc_hd__a31o_1 c653 (.A1(net317),
    .A2(net545),
    .A3(net881),
    .B1(net715),
    .X(net564));
 sky130_fd_sc_hd__sedfxtp_1 c654 (.CLK(clknet_leaf_30_clk),
    .D(net444),
    .DE(net892),
    .SCD(net563),
    .SCE(net995),
    .Q(net565));
 sky130_fd_sc_hd__a21bo_1 c655 (.A1(net69),
    .A2(net772),
    .B1_N(net700),
    .X(net566));
 sky130_fd_sc_hd__sdfxbp_1 c656 (.CLK(clknet_leaf_29_clk),
    .D(net432),
    .SCD(net881),
    .SCE(net550),
    .Q(net568),
    .Q_N(net567));
 sky130_fd_sc_hd__sedfxtp_2 c657 (.CLK(clknet_leaf_30_clk),
    .D(net564),
    .DE(net444),
    .SCD(net550),
    .SCE(net986),
    .Q(net569));
 sky130_fd_sc_hd__sedfxtp_4 c658 (.CLK(clknet_leaf_29_clk),
    .D(net563),
    .DE(net569),
    .SCD(net552),
    .SCE(net881),
    .Q(net570));
 sky130_fd_sc_hd__a21bo_2 c659 (.A1(net569),
    .A2(net570),
    .B1_N(net567),
    .X(net571));
 sky130_fd_sc_hd__xnor2_4 c66 (.A(net810),
    .B(net901),
    .Y(net4));
 sky130_fd_sc_hd__a31o_1 c660 (.A1(net339),
    .A2(net566),
    .A3(net571),
    .B1(net697),
    .X(net572));
 sky130_fd_sc_hd__sdfrbp_1 c661 (.CLK(clknet_leaf_30_clk),
    .D(net962),
    .RESET_B(net555),
    .SCD(net548),
    .SCE(net339),
    .Q(net574),
    .Q_N(net573));
 sky130_fd_sc_hd__mux4_1 c662 (.A0(net552),
    .A1(net789),
    .A2(net568),
    .A3(net563),
    .S0(net571),
    .S1(net551),
    .X(net575));
 sky130_fd_sc_hd__a41o_1 c663 (.A1(net572),
    .A2(net920),
    .A3(net570),
    .A4(net892),
    .B1(clknet_1_0__leaf_net716),
    .X(net576));
 sky130_fd_sc_hd__mux4_2 c664 (.A0(net574),
    .A1(net69),
    .A2(clknet_1_0__leaf_net576),
    .A3(net317),
    .S0(net571),
    .S1(net570),
    .X(net577));
 sky130_fd_sc_hd__sdfbbp_1 c665 (.CLK(clknet_leaf_30_clk),
    .D(net890),
    .RESET_B(clknet_1_0__leaf_net576),
    .SCD(net550),
    .SCE(net571),
    .SET_B(net573),
    .Q(net578));
 sky130_fd_sc_hd__a31o_1 c666 (.A1(net578),
    .A2(net570),
    .A3(net715),
    .B1(clknet_1_0__leaf_net716),
    .X(net579));
 sky130_fd_sc_hd__mux4_1 c667 (.A0(net348),
    .A1(net574),
    .A2(clknet_1_0__leaf_net577),
    .A3(net569),
    .S0(net563),
    .S1(clknet_1_0__leaf_net716),
    .X(net580));
 sky130_fd_sc_hd__sdfrbp_1 c668 (.CLK(clknet_leaf_29_clk),
    .D(net961),
    .RESET_B(net552),
    .SCD(net571),
    .SCE(net455),
    .Q(net581));
 sky130_fd_sc_hd__mux4_1 c669 (.A0(net579),
    .A1(net465),
    .A2(clknet_1_0__leaf_net580),
    .A3(net570),
    .S0(net569),
    .S1(net1001),
    .X(net582));
 sky130_fd_sc_hd__xnor2_1 c67 (.A(net2),
    .B(net909),
    .Y(net5));
 sky130_fd_sc_hd__mux4_1 c670 (.A0(net227),
    .A1(net574),
    .A2(clknet_1_0__leaf_net580),
    .A3(net567),
    .S0(net921),
    .S1(net717),
    .X(net583));
 sky130_fd_sc_hd__mux4_1 c671 (.A0(net581),
    .A1(net571),
    .A2(net922),
    .A3(net573),
    .S0(clknet_1_1__leaf_net580),
    .S1(net718),
    .X(net584));
 sky130_fd_sc_hd__mux4_1 c672 (.A0(net455),
    .A1(net547),
    .A2(clknet_1_0__leaf_net577),
    .A3(net482),
    .S0(net233),
    .S1(clknet_1_0__leaf_net580),
    .X(net585));
 sky130_fd_sc_hd__sdfrtn_1 c673 (.CLK_N(clknet_leaf_34_clk),
    .D(net547),
    .RESET_B(net558),
    .SCD(net772),
    .SCE(net895),
    .Q(net586));
 sky130_fd_sc_hd__a31o_1 c674 (.A1(net571),
    .A2(net545),
    .A3(net553),
    .B1(net900),
    .X(net587));
 sky130_fd_sc_hd__mux4_1 c675 (.A0(net555),
    .A1(net474),
    .A2(net895),
    .A3(net233),
    .S0(net558),
    .S1(net653),
    .X(net588));
 sky130_fd_sc_hd__sdfrtp_4 c676 (.CLK(clknet_leaf_28_clk),
    .D(net558),
    .RESET_B(clknet_1_1__leaf_net580),
    .SCD(net895),
    .SCE(net721),
    .Q(net589));
 sky130_fd_sc_hd__buf_1 c677 (.A(net759),
    .X(net590));
 sky130_fd_sc_hd__buf_1 c678 (.A(net759),
    .X(net591));
 sky130_fd_sc_hd__mux4_1 c679 (.A0(clknet_1_1__leaf_net580),
    .A1(net587),
    .A2(net895),
    .A3(net886),
    .S0(net881),
    .S1(net720),
    .X(net592));
 sky130_fd_sc_hd__a31o_1 c68 (.A1(net772),
    .A2(net901),
    .A3(net797),
    .B1(net801),
    .X(net6));
 sky130_fd_sc_hd__a21bo_1 c680 (.A1(net772),
    .A2(net789),
    .B1_N(net721),
    .X(net593));
 sky130_fd_sc_hd__a21bo_1 c681 (.A1(net545),
    .A2(net482),
    .B1_N(net589),
    .X(net594));
 sky130_fd_sc_hd__mux4_1 c682 (.A0(net558),
    .A1(net594),
    .A2(net793),
    .A3(net698),
    .S0(clknet_1_0__leaf_net716),
    .S1(net723),
    .X(net595));
 sky130_fd_sc_hd__sdfrtp_1 c683 (.CLK(clknet_leaf_25_clk),
    .D(net590),
    .RESET_B(net475),
    .SCD(net932),
    .SCE(net589),
    .Q(net596));
 sky130_fd_sc_hd__mux4_1 c684 (.A0(net475),
    .A1(net596),
    .A2(net895),
    .A3(net548),
    .S0(net589),
    .S1(net723),
    .X(net597));
 sky130_fd_sc_hd__mux4_2 c685 (.A0(net933),
    .A1(net482),
    .A2(net590),
    .A3(net596),
    .S0(clknet_1_0__leaf_net577),
    .S1(net558),
    .X(net598));
 sky130_fd_sc_hd__mux4_1 c686 (.A0(net595),
    .A1(net596),
    .A2(net558),
    .A3(net589),
    .S0(net591),
    .S1(net719),
    .X(net599));
 sky130_fd_sc_hd__sdfxtp_1 c687 (.CLK(clknet_leaf_28_clk),
    .D(net599),
    .SCD(net979),
    .SCE(net725),
    .Q(net600));
 sky130_fd_sc_hd__a31o_2 c688 (.A1(net793),
    .A2(net596),
    .A3(net589),
    .B1(net725),
    .X(net601));
 sky130_fd_sc_hd__mux4_2 c689 (.A0(net443),
    .A1(net594),
    .A2(net601),
    .A3(net593),
    .S0(net932),
    .S1(net722),
    .X(net602));
 sky130_fd_sc_hd__a21bo_4 c69 (.A1(net5),
    .A2(net901),
    .B1_N(net2),
    .X(net7));
 sky130_fd_sc_hd__a41o_1 c690 (.A1(net600),
    .A2(net594),
    .A3(net553),
    .A4(net700),
    .B1(net725),
    .X(net603));
 sky130_fd_sc_hd__a41o_1 c691 (.A1(net553),
    .A2(net603),
    .A3(net590),
    .A4(net589),
    .B1(net601),
    .X(net604));
 sky130_fd_sc_hd__sdfbbn_1 c692 (.CLK_N(clknet_leaf_25_clk),
    .D(net604),
    .RESET_B(net591),
    .SCD(net233),
    .SCE(net601),
    .SET_B(net722),
    .Q(net606),
    .Q_N(net605));
 sky130_fd_sc_hd__mux4_1 c693 (.A0(net566),
    .A1(clknet_1_1__leaf_net576),
    .A2(net475),
    .A3(net908),
    .S0(net878),
    .S1(clknet_1_1__leaf_net281),
    .X(net607));
 sky130_fd_sc_hd__mux4_1 c694 (.A0(net878),
    .A1(net548),
    .A2(net474),
    .A3(net372),
    .S0(net880),
    .S1(net722),
    .X(net608));
 sky130_fd_sc_hd__mux4_1 c695 (.A0(net550),
    .A1(net566),
    .A2(clknet_1_1__leaf_net576),
    .A3(net886),
    .S0(net878),
    .S1(net727),
    .X(net609));
 sky130_fd_sc_hd__mux4_1 c696 (.A0(net593),
    .A1(net475),
    .A2(net500),
    .A3(net878),
    .S0(clknet_1_1__leaf_net577),
    .S1(net723),
    .X(net610));
 sky130_fd_sc_hd__mux4_1 c697 (.A0(net886),
    .A1(net908),
    .A2(net779),
    .A3(net590),
    .S0(net550),
    .S1(net723),
    .X(net611));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(net590),
    .A1(net772),
    .A2(net770),
    .A3(clknet_1_0__leaf_net576),
    .S0(clknet_1_0__leaf_net716),
    .S1(net729),
    .X(net612));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(clknet_1_1__leaf_net576),
    .A1(net593),
    .A2(net500),
    .A3(clknet_1_1__leaf_net716),
    .S0(net726),
    .S1(net728),
    .X(net613));
 sky130_fd_sc_hd__xnor2_4 c70 (.A(net817),
    .B(net7),
    .Y(net8));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net589),
    .A1(net895),
    .A2(net772),
    .A3(net878),
    .S0(clknet_1_1__leaf_net577),
    .S1(net474),
    .X(net614));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(net3),
    .A1(net500),
    .A2(net878),
    .A3(net593),
    .S0(net566),
    .S1(net899),
    .X(net615));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net21),
    .A1(net589),
    .A2(net372),
    .A3(clknet_1_1__leaf_net577),
    .S0(net880),
    .S1(net730),
    .X(net616));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(clknet_1_1__leaf_net281),
    .A1(net550),
    .A2(net601),
    .A3(net605),
    .S0(net724),
    .S1(net899),
    .X(net617));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net474),
    .A1(net613),
    .A2(clknet_1_0__leaf_net598),
    .A3(net593),
    .S0(net728),
    .S1(net899),
    .X(net618));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(clknet_1_1__leaf_net386),
    .A1(net880),
    .A2(clknet_1_1__leaf_net576),
    .A3(net731),
    .S0(net732),
    .S1(net734),
    .X(net619));
 sky130_fd_sc_hd__mux4_1 c706 (.A0(clknet_1_1__leaf_net281),
    .A1(net233),
    .A2(net566),
    .A3(net727),
    .S0(net899),
    .S1(clknet_1_0__leaf_net735),
    .X(net620));
 sky130_fd_sc_hd__mux4_1 c707 (.A0(net279),
    .A1(net548),
    .A2(net895),
    .A3(net566),
    .S0(net906),
    .S1(net737),
    .X(net621));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(net878),
    .A1(net879),
    .A2(net728),
    .A3(net899),
    .S0(net733),
    .S1(net738),
    .X(net622));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(clknet_1_1__leaf_net577),
    .A1(net500),
    .A2(net601),
    .A3(net878),
    .S0(clknet_1_1__leaf_net386),
    .S1(net731),
    .X(net623));
 sky130_fd_sc_hd__xnor2_4 c71 (.A(net4),
    .B(net901),
    .Y(net9));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net491),
    .A1(net550),
    .A2(net815),
    .A3(net601),
    .S0(clknet_1_0__leaf_net736),
    .S1(net739),
    .X(net624));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net550),
    .A1(net602),
    .A2(net899),
    .A3(clknet_1_1__leaf_net735),
    .S0(net740),
    .S1(net741),
    .X(net625));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net612),
    .A1(net500),
    .A2(net731),
    .A3(net740),
    .S0(net741),
    .S1(net742),
    .X(net626));
 sky130_fd_sc_hd__mux4_1 c713 (.A0(net626),
    .A1(net886),
    .A2(net475),
    .A3(net733),
    .S0(net741),
    .S1(net742),
    .X(net627));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(clknet_1_0__leaf_net598),
    .A1(net523),
    .A2(net882),
    .A3(net880),
    .S0(net906),
    .S1(net743),
    .X(net628));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net881),
    .A1(net526),
    .A2(net886),
    .A3(net522),
    .S0(net743),
    .S1(net990),
    .X(net629));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net886),
    .A1(net233),
    .A2(net770),
    .A3(net779),
    .S0(clknet_1_1__leaf_net716),
    .S1(net899),
    .X(net630));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net465),
    .A1(net298),
    .A2(clknet_1_1__leaf_net386),
    .A3(net526),
    .S0(net886),
    .S1(net747),
    .X(net631));
 sky130_fd_sc_hd__mux4_2 c718 (.A0(net815),
    .A1(net9),
    .A2(clknet_1_1__leaf_net598),
    .A3(net886),
    .S0(clknet_1_0__leaf_net736),
    .S1(net746),
    .X(net632));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(clknet_1_1__leaf_net386),
    .A1(net606),
    .A2(net523),
    .A3(net822),
    .S0(net602),
    .S1(net746),
    .X(net633));
 sky130_fd_sc_hd__a31o_1 c72 (.A1(net8),
    .A2(net7),
    .A3(net897),
    .B1(net813),
    .X(net10));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net539),
    .A1(clknet_1_0__leaf_net632),
    .A2(net601),
    .A3(net9),
    .S0(clknet_1_1__leaf_net672),
    .S1(net746),
    .X(net634));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net879),
    .A1(clknet_1_0__leaf_net633),
    .A2(net233),
    .A3(clknet_1_1__leaf_net736),
    .S0(net743),
    .S1(net990),
    .X(net635));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net298),
    .A1(net535),
    .A2(net515),
    .A3(net601),
    .S0(clknet_1_1__leaf_net386),
    .S1(net990),
    .X(net636));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net601),
    .A1(net602),
    .A2(net372),
    .A3(net822),
    .S0(net539),
    .S1(clknet_1_1__leaf_net716),
    .X(net637));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net535),
    .A1(net464),
    .A2(net653),
    .A3(clknet_1_1__leaf_net716),
    .S0(net743),
    .S1(net746),
    .X(net638));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net372),
    .A1(net634),
    .A2(net770),
    .A3(net9),
    .S0(net747),
    .S1(net749),
    .X(net639));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net526),
    .A1(net602),
    .A2(net923),
    .A3(net233),
    .S0(net745),
    .S1(net747),
    .X(net640));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net602),
    .A1(net882),
    .A2(net526),
    .A3(net899),
    .S0(net746),
    .S1(net973),
    .X(net641));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net515),
    .A1(clknet_1_0__leaf_net632),
    .A2(net822),
    .A3(net526),
    .S0(net743),
    .S1(net748),
    .X(net642));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(net637),
    .A1(net882),
    .A2(net605),
    .A3(clknet_1_1__leaf_net672),
    .S0(net899),
    .S1(net743),
    .X(net643));
 sky130_fd_sc_hd__xnor2_4 c73 (.A(net8),
    .B(net801),
    .Y(net11));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net880),
    .A1(net606),
    .A2(net514),
    .A3(clknet_1_1__leaf_net633),
    .S0(net711),
    .S1(net751),
    .X(net644));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net606),
    .A1(clknet_1_0__leaf_net633),
    .A2(clknet_1_1__leaf_net716),
    .A3(net899),
    .S0(net746),
    .S1(net749),
    .X(net645));
 sky130_fd_sc_hd__mux4_2 c732 (.A0(clknet_1_1__leaf_net386),
    .A1(clknet_1_1__leaf_net632),
    .A2(net747),
    .A3(net752),
    .S0(net754),
    .S1(net755),
    .X(net646));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(clknet_1_1__leaf_net646),
    .A1(net880),
    .A2(net882),
    .A3(net747),
    .S0(net756),
    .S1(net757),
    .X(net647));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(clknet_1_1__leaf_net633),
    .A1(net638),
    .A2(clknet_1_0__leaf_net646),
    .A3(net747),
    .S0(net753),
    .S1(net758),
    .X(net648));
 sky130_fd_sc_hd__xnor2_4 c74 (.A(net897),
    .B(net7),
    .Y(net12));
 sky130_fd_sc_hd__a21bo_4 c75 (.A1(net10),
    .A2(net897),
    .B1_N(net901),
    .X(net13));
 sky130_fd_sc_hd__xnor2_1 c76 (.A(net12),
    .B(net897),
    .Y(net14));
 sky130_fd_sc_hd__xnor2_1 c77 (.A(net10),
    .B(net13),
    .Y(net15));
 sky130_fd_sc_hd__a41o_2 c78 (.A1(net15),
    .A2(net13),
    .A3(net5),
    .A4(net901),
    .B1(net820),
    .X(net16));
 sky130_fd_sc_hd__xnor2_2 c79 (.A(net13),
    .B(net11),
    .Y(net17));
 sky130_fd_sc_hd__a41o_1 c80 (.A1(net16),
    .A2(net818),
    .A3(net15),
    .A4(net798),
    .B1(net12),
    .X(net18));
 sky130_fd_sc_hd__a41o_4 c81 (.A1(net806),
    .A2(net7),
    .A3(net762),
    .A4(net14),
    .B1(net4),
    .X(net19));
 sky130_fd_sc_hd__xnor2_1 c82 (.A(net19),
    .B(net17),
    .Y(net20));
 sky130_fd_sc_hd__mux4_2 c83 (.A0(net14),
    .A1(net7),
    .A2(net20),
    .A3(net19),
    .S0(net16),
    .S1(net13),
    .X(net21));
 sky130_fd_sc_hd__xnor2_4 c84 (.A(net801),
    .B(net2),
    .Y(net22));
 sky130_fd_sc_hd__a21bo_4 c85 (.A1(net19),
    .A2(net761),
    .B1_N(net16),
    .X(net23));
 sky130_fd_sc_hd__xnor2_2 c86 (.A(net16),
    .B(net22),
    .Y(net24));
 sky130_fd_sc_hd__a31o_4 c87 (.A1(net24),
    .A2(net2),
    .A3(net22),
    .B1(net19),
    .X(net25));
 sky130_fd_sc_hd__xnor2_1 c88 (.A(net814),
    .B(net11),
    .Y(net26));
 sky130_fd_sc_hd__a21bo_2 c89 (.A1(net26),
    .A2(net797),
    .B1_N(net24),
    .X(net27));
 sky130_fd_sc_hd__xnor2_4 c90 (.A(net25),
    .B(net23),
    .Y(net28));
 sky130_fd_sc_hd__a31o_1 c91 (.A1(net2),
    .A2(net23),
    .A3(net28),
    .B1(net4),
    .X(net29));
 sky130_fd_sc_hd__xnor2_2 c92 (.A(net762),
    .B(net22),
    .Y(net30));
 sky130_fd_sc_hd__xnor2_4 c93 (.A(net25),
    .B(net888),
    .Y(net31));
 sky130_fd_sc_hd__a31o_1 c94 (.A1(net30),
    .A2(net4),
    .A3(net24),
    .B1(net797),
    .X(net32));
 sky130_fd_sc_hd__a31o_1 c95 (.A1(net32),
    .A2(net16),
    .A3(net23),
    .B1(net26),
    .X(net33));
 sky130_fd_sc_hd__a31o_1 c96 (.A1(net32),
    .A2(net31),
    .A3(net27),
    .B1(net16),
    .X(net34));
 sky130_fd_sc_hd__a31o_1 c97 (.A1(net26),
    .A2(net19),
    .A3(net803),
    .B1(net11),
    .X(net35));
 sky130_fd_sc_hd__xnor2_2 c98 (.A(net23),
    .B(net28),
    .Y(net36));
 sky130_fd_sc_hd__a21bo_1 c99 (.A1(net33),
    .A2(net32),
    .B1_N(net31),
    .X(net37));
 sky130_fd_sc_hd__mux4_1 merge740 (.A0(net570),
    .A1(net589),
    .A2(net547),
    .A3(net586),
    .S0(net474),
    .S1(net699),
    .X(net649));
 sky130_fd_sc_hd__dfxbp_1 s741 (.CLK(clknet_leaf_7_clk),
    .D(net39),
    .Q(net651),
    .Q_N(net650));
 sky130_fd_sc_hd__dfxbp_2 s742 (.CLK(clknet_leaf_7_clk),
    .D(net41),
    .Q(net867),
    .Q_N(net652));
 sky130_fd_sc_hd__dfxtp_1 s743 (.CLK(clknet_leaf_8_clk),
    .D(net65),
    .Q(net854));
 sky130_fd_sc_hd__dfxtp_1 s744 (.CLK(clknet_leaf_9_clk),
    .D(net66),
    .Q(net847));
 sky130_fd_sc_hd__dfxtp_2 s745 (.CLK(clknet_leaf_0_clk),
    .D(net126),
    .Q(net653));
 sky130_fd_sc_hd__dlclkp_1 s746 (.CLK(clknet_leaf_0_clk),
    .GATE(net129),
    .GCLK(net859));
 sky130_fd_sc_hd__dlclkp_2 s747 (.CLK(clknet_leaf_0_clk),
    .GATE(net146),
    .GCLK(net654));
 sky130_fd_sc_hd__dlclkp_4 s748 (.CLK(clknet_leaf_5_clk),
    .GATE(net152),
    .GCLK(net655));
 sky130_fd_sc_hd__dlxbn_1 s749 (.D(net153),
    .GATE_N(clknet_leaf_4_clk),
    .Q(net657),
    .Q_N(net656));
 sky130_fd_sc_hd__dlxbn_1 s750 (.D(net177),
    .GATE_N(clknet_leaf_13_clk),
    .Q(net659),
    .Q_N(net658));
 sky130_fd_sc_hd__dlxbp_1 s751 (.D(net178),
    .GATE(clknet_leaf_10_clk),
    .Q(net869),
    .Q_N(net660));
 sky130_fd_sc_hd__dlxtn_2 s752 (.D(net179),
    .GATE_N(clknet_leaf_10_clk),
    .Q(net875));
 sky130_fd_sc_hd__dlxtn_1 s753 (.D(net189),
    .GATE_N(clknet_leaf_9_clk),
    .Q(net661));
 sky130_fd_sc_hd__dlxtn_1 s754 (.D(net197),
    .GATE_N(clknet_leaf_10_clk),
    .Q(net828));
 sky130_fd_sc_hd__dlxtp_1 s755 (.D(net218),
    .GATE(clknet_leaf_41_clk),
    .Q(net662));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s756 (.D(net261),
    .SLEEP_B(clknet_leaf_1_clk),
    .Q(net663));
 sky130_fd_sc_hd__dfxbp_1 s757 (.CLK(clknet_leaf_2_clk),
    .D(net269),
    .Q(net665),
    .Q_N(net664));
 sky130_fd_sc_hd__dfxbp_1 s758 (.CLK(clknet_leaf_3_clk),
    .D(net278),
    .Q(net667),
    .Q_N(net666));
 sky130_fd_sc_hd__dfxtp_1 s759 (.CLK(clknet_leaf_4_clk),
    .D(net284),
    .Q(net668));
 sky130_fd_sc_hd__dfxtp_1 s760 (.CLK(clknet_leaf_3_clk),
    .D(net285),
    .Q(net669));
 sky130_fd_sc_hd__dfxtp_1 s761 (.CLK(clknet_leaf_4_clk),
    .D(net294),
    .Q(net670));
 sky130_fd_sc_hd__dlclkp_1 s762 (.CLK(clknet_leaf_12_clk),
    .GATE(net302),
    .GCLK(net671));
 sky130_fd_sc_hd__dlclkp_2 s763 (.CLK(clknet_leaf_12_clk),
    .GATE(net305),
    .GCLK(net672));
 sky130_fd_sc_hd__dlclkp_4 s764 (.CLK(clknet_leaf_11_clk),
    .GATE(net306),
    .GCLK(net868));
 sky130_fd_sc_hd__dlxbn_1 s765 (.D(net307),
    .GATE_N(clknet_leaf_11_clk),
    .Q(net870),
    .Q_N(net865));
 sky130_fd_sc_hd__dlxbn_1 s766 (.D(net308),
    .GATE_N(clknet_leaf_11_clk),
    .Q(net866),
    .Q_N(net673));
 sky130_fd_sc_hd__dlxbp_1 s767 (.D(net309),
    .GATE(clknet_leaf_11_clk),
    .Q(net864),
    .Q_N(net674));
 sky130_fd_sc_hd__dlxtn_4 s768 (.D(net329),
    .GATE_N(clknet_leaf_40_clk),
    .Q(net675));
 sky130_fd_sc_hd__dlxtn_1 s769 (.D(net331),
    .GATE_N(clknet_leaf_40_clk),
    .Q(net676));
 sky130_fd_sc_hd__dlxtn_1 s770 (.D(net334),
    .GATE_N(clknet_leaf_33_clk),
    .Q(net677));
 sky130_fd_sc_hd__dlxtp_1 s771 (.D(net341),
    .GATE(clknet_leaf_37_clk),
    .Q(net678));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s772 (.D(net343),
    .SLEEP_B(clknet_leaf_37_clk),
    .Q(net679));
 sky130_fd_sc_hd__dfxbp_1 s773 (.CLK(clknet_leaf_37_clk),
    .D(net357),
    .Q(net680));
 sky130_fd_sc_hd__dfxbp_1 s774 (.CLK(clknet_leaf_37_clk),
    .D(net362),
    .Q(net682),
    .Q_N(net681));
 sky130_fd_sc_hd__dfxtp_1 s775 (.CLK(clknet_leaf_37_clk),
    .D(net374),
    .Q(net683));
 sky130_fd_sc_hd__dfxtp_1 s776 (.CLK(clknet_leaf_36_clk),
    .D(net376),
    .Q(net684));
 sky130_fd_sc_hd__dfxtp_1 s777 (.CLK(clknet_leaf_35_clk),
    .D(net378),
    .Q(net685));
 sky130_fd_sc_hd__dlclkp_1 s778 (.CLK(clknet_leaf_35_clk),
    .GATE(net379),
    .GCLK(net686));
 sky130_fd_sc_hd__dlclkp_2 s779 (.CLK(clknet_leaf_2_clk),
    .GATE(net384),
    .GCLK(net687));
 sky130_fd_sc_hd__dlclkp_4 s780 (.CLK(clknet_leaf_15_clk),
    .GATE(net392),
    .GCLK(net688));
 sky130_fd_sc_hd__dlxbn_1 s781 (.D(net394),
    .GATE_N(clknet_leaf_14_clk),
    .Q(net689));
 sky130_fd_sc_hd__dlxbn_1 s782 (.D(net398),
    .GATE_N(clknet_leaf_16_clk),
    .Q(net691),
    .Q_N(net690));
 sky130_fd_sc_hd__dlxbp_1 s783 (.D(net402),
    .GATE(clknet_leaf_16_clk),
    .Q(net693),
    .Q_N(net692));
 sky130_fd_sc_hd__dlxtn_2 s784 (.D(net406),
    .GATE_N(clknet_leaf_18_clk),
    .Q(net694));
 sky130_fd_sc_hd__dlxtn_1 s785 (.D(net410),
    .GATE_N(clknet_leaf_12_clk),
    .Q(net848));
 sky130_fd_sc_hd__dlxtn_1 s786 (.D(net411),
    .GATE_N(clknet_leaf_12_clk),
    .Q(net860));
 sky130_fd_sc_hd__dlxtp_1 s787 (.D(net414),
    .GATE(clknet_leaf_14_clk),
    .Q(net695));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s788 (.D(net418),
    .SLEEP_B(clknet_leaf_17_clk),
    .Q(net858));
 sky130_fd_sc_hd__dfxbp_1 s789 (.CLK(clknet_leaf_34_clk),
    .D(net451),
    .Q(net696));
 sky130_fd_sc_hd__dfxbp_1 s790 (.CLK(clknet_leaf_34_clk),
    .D(net456),
    .Q(net698),
    .Q_N(net697));
 sky130_fd_sc_hd__dfxtp_1 s791 (.CLK(clknet_leaf_33_clk),
    .D(net460),
    .Q(net699));
 sky130_fd_sc_hd__dfxtp_1 s792 (.CLK(clknet_leaf_34_clk),
    .D(net466),
    .Q(net700));
 sky130_fd_sc_hd__dfxtp_1 s793 (.CLK(clknet_leaf_35_clk),
    .D(net481),
    .Q(net701));
 sky130_fd_sc_hd__dlclkp_1 s794 (.CLK(clknet_leaf_34_clk),
    .GATE(net486),
    .GCLK(net702));
 sky130_fd_sc_hd__dlclkp_2 s795 (.CLK(clknet_leaf_24_clk),
    .GATE(net492),
    .GCLK(net834));
 sky130_fd_sc_hd__dlclkp_4 s796 (.CLK(clknet_leaf_24_clk),
    .GATE(net499),
    .GCLK(net703));
 sky130_fd_sc_hd__dlxbn_1 s797 (.D(net504),
    .GATE_N(clknet_leaf_23_clk),
    .Q(net704));
 sky130_fd_sc_hd__dlxbn_1 s798 (.D(net507),
    .GATE_N(clknet_leaf_23_clk),
    .Q(net705));
 sky130_fd_sc_hd__dlxbp_1 s799 (.D(net510),
    .GATE(clknet_leaf_27_clk),
    .Q(net824));
 sky130_fd_sc_hd__dlxtn_1 s800 (.D(net519),
    .GATE_N(clknet_leaf_15_clk),
    .Q(net706));
 sky130_fd_sc_hd__dlxtn_1 s801 (.D(net520),
    .GATE_N(clknet_leaf_22_clk),
    .Q(net707));
 sky130_fd_sc_hd__dlxtn_2 s802 (.D(net521),
    .GATE_N(clknet_leaf_16_clk),
    .Q(net708));
 sky130_fd_sc_hd__dlxtp_1 s803 (.D(net529),
    .GATE(clknet_leaf_16_clk),
    .Q(net709));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s804 (.D(net536),
    .SLEEP_B(clknet_leaf_17_clk),
    .Q(net710));
 sky130_fd_sc_hd__dfxbp_1 s805 (.CLK(clknet_leaf_19_clk),
    .D(net537),
    .Q(net711));
 sky130_fd_sc_hd__dfxbp_1 s806 (.CLK(clknet_leaf_19_clk),
    .D(net538),
    .Q(net712));
 sky130_fd_sc_hd__dfxtp_1 s807 (.CLK(clknet_leaf_31_clk),
    .D(net554),
    .Q(net713));
 sky130_fd_sc_hd__dfxtp_1 s808 (.CLK(clknet_leaf_30_clk),
    .D(net560),
    .Q(net714));
 sky130_fd_sc_hd__dfxtp_1 s809 (.CLK(clknet_leaf_30_clk),
    .D(net561),
    .Q(net715));
 sky130_fd_sc_hd__dlclkp_1 s810 (.CLK(clknet_leaf_29_clk),
    .GATE(net575),
    .GCLK(net716));
 sky130_fd_sc_hd__dlclkp_2 s811 (.CLK(clknet_leaf_29_clk),
    .GATE(net582),
    .GCLK(net717));
 sky130_fd_sc_hd__dlclkp_4 s812 (.CLK(clknet_leaf_28_clk),
    .GATE(net583),
    .GCLK(net718));
 sky130_fd_sc_hd__dlxbn_1 s813 (.D(net584),
    .GATE_N(clknet_leaf_28_clk),
    .Q(net719));
 sky130_fd_sc_hd__dlxbn_1 s814 (.D(net585),
    .GATE_N(clknet_leaf_28_clk),
    .Q(net721),
    .Q_N(net720));
 sky130_fd_sc_hd__dlxbp_1 s815 (.D(net588),
    .GATE(clknet_leaf_25_clk),
    .Q(net723),
    .Q_N(net722));
 sky130_fd_sc_hd__dlxtn_1 s816 (.D(net592),
    .GATE_N(clknet_leaf_28_clk),
    .Q(net724));
 sky130_fd_sc_hd__dlxtn_1 s817 (.D(net597),
    .GATE_N(clknet_leaf_28_clk),
    .Q(net725));
 sky130_fd_sc_hd__dlxtn_1 s818 (.D(net607),
    .GATE_N(clknet_leaf_25_clk),
    .Q(net726));
 sky130_fd_sc_hd__dlxtp_1 s819 (.D(net608),
    .GATE(clknet_leaf_25_clk),
    .Q(net727));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s820 (.D(net609),
    .SLEEP_B(clknet_leaf_25_clk),
    .Q(net728));
 sky130_fd_sc_hd__dfxbp_1 s821 (.CLK(clknet_leaf_27_clk),
    .D(net610),
    .Q(net729));
 sky130_fd_sc_hd__dfxbp_1 s822 (.CLK(clknet_leaf_27_clk),
    .D(net611),
    .Q(net730));
 sky130_fd_sc_hd__dfxtp_1 s823 (.CLK(clknet_leaf_25_clk),
    .D(net614),
    .Q(net731));
 sky130_fd_sc_hd__dfxtp_1 s824 (.CLK(clknet_leaf_26_clk),
    .D(net615),
    .Q(net732));
 sky130_fd_sc_hd__dfxtp_1 s825 (.CLK(clknet_leaf_27_clk),
    .D(net616),
    .Q(net733));
 sky130_fd_sc_hd__dlclkp_1 s826 (.CLK(clknet_leaf_26_clk),
    .GATE(net617),
    .GCLK(net734));
 sky130_fd_sc_hd__dlclkp_2 s827 (.CLK(clknet_leaf_26_clk),
    .GATE(net618),
    .GCLK(net735));
 sky130_fd_sc_hd__dlclkp_4 s828 (.CLK(clknet_leaf_21_clk),
    .GATE(net619),
    .GCLK(net736));
 sky130_fd_sc_hd__dlxbn_1 s829 (.D(net620),
    .GATE_N(clknet_leaf_25_clk),
    .Q(net737));
 sky130_fd_sc_hd__dlxbn_1 s830 (.D(net621),
    .GATE_N(clknet_leaf_26_clk),
    .Q(net738));
 sky130_fd_sc_hd__dlxbp_1 s831 (.D(net622),
    .GATE(clknet_leaf_26_clk),
    .Q(net739));
 sky130_fd_sc_hd__dlxtn_1 s832 (.D(net623),
    .GATE_N(clknet_leaf_26_clk),
    .Q(net740));
 sky130_fd_sc_hd__dlxtn_1 s833 (.D(net624),
    .GATE_N(clknet_leaf_26_clk),
    .Q(net741));
 sky130_fd_sc_hd__dlxtn_1 s834 (.D(net625),
    .GATE_N(clknet_leaf_27_clk),
    .Q(net742));
 sky130_fd_sc_hd__dlxtp_1 s835 (.D(net627),
    .GATE(clknet_leaf_21_clk),
    .Q(net743));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s836 (.D(net628),
    .SLEEP_B(clknet_leaf_22_clk),
    .Q(net744));
 sky130_fd_sc_hd__dfxbp_1 s837 (.CLK(clknet_leaf_23_clk),
    .D(net629),
    .Q(net745));
 sky130_fd_sc_hd__dfxbp_2 s838 (.CLK(clknet_leaf_20_clk),
    .D(net630),
    .Q(net747),
    .Q_N(net746));
 sky130_fd_sc_hd__dfxtp_1 s839 (.CLK(clknet_leaf_19_clk),
    .D(net631),
    .Q(net748));
 sky130_fd_sc_hd__dfxtp_1 s840 (.CLK(clknet_leaf_21_clk),
    .D(net635),
    .Q(net749));
 sky130_fd_sc_hd__dfxtp_1 s841 (.CLK(clknet_leaf_22_clk),
    .D(net636),
    .Q(net750));
 sky130_fd_sc_hd__dlclkp_1 s842 (.CLK(clknet_leaf_20_clk),
    .GATE(net639),
    .GCLK(net751));
 sky130_fd_sc_hd__dlclkp_2 s843 (.CLK(clknet_leaf_19_clk),
    .GATE(net640),
    .GCLK(net752));
 sky130_fd_sc_hd__dlclkp_4 s844 (.CLK(clknet_leaf_20_clk),
    .GATE(net641),
    .GCLK(net753));
 sky130_fd_sc_hd__dlxbn_1 s845 (.D(net642),
    .GATE_N(clknet_leaf_19_clk),
    .Q(net754));
 sky130_fd_sc_hd__dlxbn_1 s846 (.D(net643),
    .GATE_N(clknet_leaf_21_clk),
    .Q(net823));
 sky130_fd_sc_hd__dlxbp_1 s847 (.D(net644),
    .GATE(clknet_leaf_20_clk),
    .Q(net756),
    .Q_N(net755));
 sky130_fd_sc_hd__dlxtn_1 s848 (.D(net645),
    .GATE_N(clknet_leaf_20_clk),
    .Q(net757));
 sky130_fd_sc_hd__dlxtn_1 s849 (.D(net647),
    .GATE_N(clknet_leaf_20_clk),
    .Q(net758));
 sky130_fd_sc_hd__dlxtn_4 s850 (.D(net648),
    .GATE_N(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dlxtp_1 s851 (.D(net649),
    .GATE(clknet_leaf_28_clk),
    .Q(net759));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(in0),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_8 input2 (.A(in1),
    .X(net761));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(in10),
    .X(net762));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(in11),
    .X(net763));
 sky130_fd_sc_hd__buf_1 input5 (.A(in12),
    .X(net764));
 sky130_fd_sc_hd__buf_2 input6 (.A(in13),
    .X(net765));
 sky130_fd_sc_hd__buf_2 input7 (.A(in14),
    .X(net766));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(in15),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(in16),
    .X(net768));
 sky130_fd_sc_hd__buf_2 input10 (.A(in17),
    .X(net769));
 sky130_fd_sc_hd__clkbuf_8 input11 (.A(in18),
    .X(net770));
 sky130_fd_sc_hd__buf_4 input12 (.A(in19),
    .X(net771));
 sky130_fd_sc_hd__buf_4 input13 (.A(in2),
    .X(net772));
 sky130_fd_sc_hd__buf_2 input14 (.A(in20),
    .X(net773));
 sky130_fd_sc_hd__buf_1 input15 (.A(in21),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(in22),
    .X(net775));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(in23),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(in24),
    .X(net777));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(in25),
    .X(net778));
 sky130_fd_sc_hd__buf_6 input20 (.A(in26),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(in27),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(in28),
    .X(net781));
 sky130_fd_sc_hd__clkbuf_4 input23 (.A(in29),
    .X(net782));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(in3),
    .X(net783));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(in30),
    .X(net784));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(in31),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(in32),
    .X(net786));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(in33),
    .X(net787));
 sky130_fd_sc_hd__buf_1 input29 (.A(in34),
    .X(net788));
 sky130_fd_sc_hd__buf_4 input30 (.A(in35),
    .X(net789));
 sky130_fd_sc_hd__buf_1 input31 (.A(in36),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(in37),
    .X(net791));
 sky130_fd_sc_hd__buf_4 input33 (.A(in38),
    .X(net792));
 sky130_fd_sc_hd__buf_1 input34 (.A(in39),
    .X(net793));
 sky130_fd_sc_hd__buf_2 input35 (.A(in4),
    .X(net794));
 sky130_fd_sc_hd__dlymetal6s2s_1 input36 (.A(in40),
    .X(net795));
 sky130_fd_sc_hd__buf_1 input37 (.A(in41),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(in42),
    .X(net797));
 sky130_fd_sc_hd__buf_1 input39 (.A(in43),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(in44),
    .X(net799));
 sky130_fd_sc_hd__clkbuf_4 input41 (.A(in45),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(in46),
    .X(net801));
 sky130_fd_sc_hd__buf_2 input43 (.A(in47),
    .X(net802));
 sky130_fd_sc_hd__buf_2 input44 (.A(in48),
    .X(net803));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(in49),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(in5),
    .X(net805));
 sky130_fd_sc_hd__buf_1 input47 (.A(in50),
    .X(net806));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(in51),
    .X(net807));
 sky130_fd_sc_hd__buf_1 input49 (.A(in52),
    .X(net808));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(in53),
    .X(net809));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(in54),
    .X(net810));
 sky130_fd_sc_hd__dlymetal6s2s_1 input52 (.A(in55),
    .X(net811));
 sky130_fd_sc_hd__buf_1 input53 (.A(in56),
    .X(net812));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(in57),
    .X(net813));
 sky130_fd_sc_hd__buf_1 input55 (.A(in58),
    .X(net814));
 sky130_fd_sc_hd__buf_1 input56 (.A(in59),
    .X(net815));
 sky130_fd_sc_hd__buf_4 input57 (.A(in6),
    .X(net816));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(in60),
    .X(net817));
 sky130_fd_sc_hd__buf_1 input59 (.A(in61),
    .X(net818));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(in7),
    .X(net819));
 sky130_fd_sc_hd__buf_4 input61 (.A(in8),
    .X(net820));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(in9),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net822),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output64 (.A(net823),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output65 (.A(net824),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output66 (.A(net825),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(clknet_1_1__leaf_net826),
    .X(out12));
 sky130_fd_sc_hd__clkbuf_4 output68 (.A(net827),
    .X(out13));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net828),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output70 (.A(net829),
    .X(out15));
 sky130_fd_sc_hd__clkbuf_4 output71 (.A(net830),
    .X(out16));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(clknet_1_1__leaf_net831),
    .X(out17));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net832),
    .X(out18));
 sky130_fd_sc_hd__clkbuf_4 output74 (.A(net833),
    .X(out19));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(clknet_1_1__leaf_net834),
    .X(out20));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net835),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_4 output77 (.A(net836),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output78 (.A(net837),
    .X(out24));
 sky130_fd_sc_hd__clkbuf_4 output79 (.A(net838),
    .X(out25));
 sky130_fd_sc_hd__buf_2 output80 (.A(net839),
    .X(out27));
 sky130_fd_sc_hd__clkbuf_4 output81 (.A(net840),
    .X(out28));
 sky130_fd_sc_hd__clkbuf_4 output82 (.A(net841),
    .X(out29));
 sky130_fd_sc_hd__buf_2 output83 (.A(net842),
    .X(out3));
 sky130_fd_sc_hd__clkbuf_4 output84 (.A(net843),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output85 (.A(net844),
    .X(out31));
 sky130_fd_sc_hd__clkbuf_4 output86 (.A(net905),
    .X(out32));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(clknet_1_1__leaf_net846),
    .X(out33));
 sky130_fd_sc_hd__clkbuf_4 output88 (.A(net847),
    .X(out34));
 sky130_fd_sc_hd__clkbuf_4 output89 (.A(net848),
    .X(out35));
 sky130_fd_sc_hd__clkbuf_4 output90 (.A(net849),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_4 output91 (.A(net850),
    .X(out37));
 sky130_fd_sc_hd__clkbuf_4 output92 (.A(net851),
    .X(out38));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net852),
    .X(out39));
 sky130_fd_sc_hd__clkbuf_4 output94 (.A(net853),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_4 output95 (.A(net854),
    .X(out40));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(clknet_1_1__leaf_net855),
    .X(out41));
 sky130_fd_sc_hd__clkbuf_1 output97 (.A(net856),
    .X(out42));
 sky130_fd_sc_hd__clkbuf_4 output98 (.A(net857),
    .X(out43));
 sky130_fd_sc_hd__clkbuf_4 output99 (.A(net858),
    .X(out44));
 sky130_fd_sc_hd__clkbuf_1 output100 (.A(clknet_1_1__leaf_net859),
    .X(out45));
 sky130_fd_sc_hd__clkbuf_4 output101 (.A(net860),
    .X(out46));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(net861),
    .X(out47));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net862),
    .X(out48));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net863),
    .X(out49));
 sky130_fd_sc_hd__clkbuf_4 output105 (.A(net864),
    .X(out50));
 sky130_fd_sc_hd__clkbuf_4 output106 (.A(net865),
    .X(out51));
 sky130_fd_sc_hd__clkbuf_4 output107 (.A(net866),
    .X(out52));
 sky130_fd_sc_hd__clkbuf_4 output108 (.A(net867),
    .X(out53));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(net868),
    .X(out55));
 sky130_fd_sc_hd__clkbuf_4 output110 (.A(net869),
    .X(out56));
 sky130_fd_sc_hd__clkbuf_4 output111 (.A(net870),
    .X(out57));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(clknet_1_1__leaf_net871),
    .X(out58));
 sky130_fd_sc_hd__clkbuf_4 output113 (.A(net872),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output114 (.A(net873),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(clknet_1_1__leaf_net874),
    .X(out61));
 sky130_fd_sc_hd__clkbuf_4 output116 (.A(net875),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output117 (.A(net876),
    .X(out8));
 sky130_fd_sc_hd__clkbuf_4 output118 (.A(net877),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_4 fanout119 (.A(net491),
    .X(net878));
 sky130_fd_sc_hd__buf_4 max_cap120 (.A(net444),
    .X(net879));
 sky130_fd_sc_hd__buf_4 fanout121 (.A(net842),
    .X(net880));
 sky130_fd_sc_hd__buf_4 fanout122 (.A(net440),
    .X(net881));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout123 (.A(net440),
    .X(net882));
 sky130_fd_sc_hd__buf_4 max_cap124 (.A(net310),
    .X(net883));
 sky130_fd_sc_hd__buf_4 fanout125 (.A(net138),
    .X(net884));
 sky130_fd_sc_hd__clkbuf_8 fanout126 (.A(net211),
    .X(net885));
 sky130_fd_sc_hd__buf_2 fanout127 (.A(net929),
    .X(net886));
 sky130_fd_sc_hd__buf_4 fanout128 (.A(net102),
    .X(net887));
 sky130_fd_sc_hd__buf_4 max_cap129 (.A(net24),
    .X(net888));
 sky130_fd_sc_hd__buf_4 max_cap130 (.A(net423),
    .X(net889));
 sky130_fd_sc_hd__buf_4 max_cap131 (.A(net202),
    .X(net890));
 sky130_fd_sc_hd__clkbuf_4 fanout132 (.A(net892),
    .X(net891));
 sky130_fd_sc_hd__buf_2 fanout133 (.A(net422),
    .X(net892));
 sky130_fd_sc_hd__buf_12 fanout134 (.A(net199),
    .X(net893));
 sky130_fd_sc_hd__buf_4 fanout135 (.A(net314),
    .X(net894));
 sky130_fd_sc_hd__clkbuf_4 fanout136 (.A(net314),
    .X(net895));
 sky130_fd_sc_hd__buf_4 max_cap137 (.A(net83),
    .X(net896));
 sky130_fd_sc_hd__buf_4 fanout138 (.A(net9),
    .X(net897));
 sky130_fd_sc_hd__clkbuf_4 fanout139 (.A(net140),
    .X(net898));
 sky130_fd_sc_hd__clkbuf_4 fanout140 (.A(net731),
    .X(net899));
 sky130_fd_sc_hd__buf_4 fanout141 (.A(net653),
    .X(net900));
 sky130_fd_sc_hd__clkbuf_8 fanout142 (.A(net3),
    .X(net901));
 sky130_fd_sc_hd__buf_2 fanout143 (.A(net904),
    .X(net902));
 sky130_fd_sc_hd__clkbuf_2 fanout144 (.A(net904),
    .X(net903));
 sky130_fd_sc_hd__buf_2 fanout145 (.A(net905),
    .X(net904));
 sky130_fd_sc_hd__buf_2 fanout146 (.A(net845),
    .X(net905));
 sky130_fd_sc_hd__buf_12 fanout147 (.A(net70),
    .X(net906));
 sky130_fd_sc_hd__clkbuf_8 fanout148 (.A(net857),
    .X(net907));
 sky130_fd_sc_hd__clkbuf_4 fanout149 (.A(net815),
    .X(net908));
 sky130_fd_sc_hd__buf_4 fanout150 (.A(net807),
    .X(net909));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_36_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_37_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_38_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_40_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_41_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_42_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_43_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net646 (.A(net646),
    .X(clknet_0_net646));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net646 (.A(clknet_0_net646),
    .X(clknet_1_0__leaf_net646));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net646 (.A(clknet_0_net646),
    .X(clknet_1_1__leaf_net646));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net736 (.A(net736),
    .X(clknet_0_net736));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net736 (.A(clknet_0_net736),
    .X(clknet_1_0__leaf_net736));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net736 (.A(clknet_0_net736),
    .X(clknet_1_1__leaf_net736));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net632 (.A(net632),
    .X(clknet_0_net632));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net632 (.A(clknet_0_net632),
    .X(clknet_1_0__leaf_net632));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net632 (.A(clknet_0_net632),
    .X(clknet_1_1__leaf_net632));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net735 (.A(net735),
    .X(clknet_0_net735));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net735 (.A(clknet_0_net735),
    .X(clknet_1_0__leaf_net735));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net735 (.A(clknet_0_net735),
    .X(clknet_1_1__leaf_net735));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net716 (.A(net716),
    .X(clknet_0_net716));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net716 (.A(clknet_0_net716),
    .X(clknet_1_0__leaf_net716));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net716 (.A(clknet_0_net716),
    .X(clknet_1_1__leaf_net716));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net580 (.A(net580),
    .X(clknet_0_net580));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net580 (.A(clknet_0_net580),
    .X(clknet_1_0__leaf_net580));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net580 (.A(clknet_0_net580),
    .X(clknet_1_1__leaf_net580));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net576 (.A(net576),
    .X(clknet_0_net576));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net576 (.A(clknet_0_net576),
    .X(clknet_1_0__leaf_net576));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net576 (.A(clknet_0_net576),
    .X(clknet_1_1__leaf_net576));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net577 (.A(net577),
    .X(clknet_0_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net577 (.A(clknet_0_net577),
    .X(clknet_1_0__leaf_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net577 (.A(clknet_0_net577),
    .X(clknet_1_1__leaf_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net598 (.A(net598),
    .X(clknet_0_net598));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net598 (.A(clknet_0_net598),
    .X(clknet_1_0__leaf_net598));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net598 (.A(clknet_0_net598),
    .X(clknet_1_1__leaf_net598));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net834 (.A(net834),
    .X(clknet_0_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net834 (.A(clknet_0_net834),
    .X(clknet_1_0__leaf_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net834 (.A(clknet_0_net834),
    .X(clknet_1_1__leaf_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net531 (.A(net531),
    .X(clknet_0_net531));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net531 (.A(clknet_0_net531),
    .X(clknet_1_0__leaf_net531));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net531 (.A(clknet_0_net531),
    .X(clknet_1_1__leaf_net531));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net702 (.A(net702),
    .X(clknet_0_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net702 (.A(clknet_0_net702),
    .X(clknet_1_0__leaf_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net702 (.A(clknet_0_net702),
    .X(clknet_1_1__leaf_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net826 (.A(net826),
    .X(clknet_0_net826));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net826 (.A(clknet_0_net826),
    .X(clknet_1_0__leaf_net826));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net826 (.A(clknet_0_net826),
    .X(clknet_1_1__leaf_net826));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net687 (.A(net687),
    .X(clknet_0_net687));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net687 (.A(clknet_0_net687),
    .X(clknet_1_0__leaf_net687));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net687 (.A(clknet_0_net687),
    .X(clknet_1_1__leaf_net687));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net846 (.A(net846),
    .X(clknet_0_net846));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net846 (.A(clknet_0_net846),
    .X(clknet_1_0__leaf_net846));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net846 (.A(clknet_0_net846),
    .X(clknet_1_1__leaf_net846));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net501 (.A(net501),
    .X(clknet_0_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net501 (.A(clknet_0_net501),
    .X(clknet_1_0__leaf_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net501 (.A(clknet_0_net501),
    .X(clknet_1_1__leaf_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net386 (.A(net386),
    .X(clknet_0_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net386 (.A(clknet_0_net386),
    .X(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net386 (.A(clknet_0_net386),
    .X(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net633 (.A(net633),
    .X(clknet_0_net633));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net633 (.A(clknet_0_net633),
    .X(clknet_1_0__leaf_net633));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net633 (.A(clknet_0_net633),
    .X(clknet_1_1__leaf_net633));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net393 (.A(net393),
    .X(clknet_0_net393));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net393 (.A(clknet_0_net393),
    .X(clknet_1_0__leaf_net393));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net393 (.A(clknet_0_net393),
    .X(clknet_1_1__leaf_net393));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net389 (.A(net389),
    .X(clknet_0_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_0__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_1__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net686 (.A(net686),
    .X(clknet_0_net686));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net686 (.A(clknet_0_net686),
    .X(clknet_1_0__leaf_net686));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net686 (.A(clknet_0_net686),
    .X(clknet_1_1__leaf_net686));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net672 (.A(net672),
    .X(clknet_0_net672));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net672 (.A(clknet_0_net672),
    .X(clknet_1_0__leaf_net672));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net672 (.A(clknet_0_net672),
    .X(clknet_1_1__leaf_net672));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net403 (.A(net403),
    .X(clknet_0_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net403 (.A(clknet_0_net403),
    .X(clknet_1_0__leaf_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net403 (.A(clknet_0_net403),
    .X(clknet_1_1__leaf_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net831 (.A(net831),
    .X(clknet_0_net831));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net831 (.A(clknet_0_net831),
    .X(clknet_1_0__leaf_net831));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net831 (.A(clknet_0_net831),
    .X(clknet_1_1__leaf_net831));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net871 (.A(net871),
    .X(clknet_0_net871));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net871 (.A(clknet_0_net871),
    .X(clknet_1_0__leaf_net871));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net871 (.A(clknet_0_net871),
    .X(clknet_1_1__leaf_net871));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net671 (.A(net671),
    .X(clknet_0_net671));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net671 (.A(clknet_0_net671),
    .X(clknet_1_0__leaf_net671));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net671 (.A(clknet_0_net671),
    .X(clknet_1_1__leaf_net671));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net655 (.A(net655),
    .X(clknet_0_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net655 (.A(clknet_0_net655),
    .X(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net655 (.A(clknet_0_net655),
    .X(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net299 (.A(net299),
    .X(clknet_0_net299));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net299 (.A(clknet_0_net299),
    .X(clknet_1_0__leaf_net299));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net299 (.A(clknet_0_net299),
    .X(clknet_1_1__leaf_net299));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net154 (.A(net154),
    .X(clknet_0_net154));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net154 (.A(clknet_0_net154),
    .X(clknet_1_0__leaf_net154));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net154 (.A(clknet_0_net154),
    .X(clknet_1_1__leaf_net154));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net275 (.A(net275),
    .X(clknet_0_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net275 (.A(clknet_0_net275),
    .X(clknet_1_0__leaf_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net275 (.A(clknet_0_net275),
    .X(clknet_1_1__leaf_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net281 (.A(net281),
    .X(clknet_0_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net281 (.A(clknet_0_net281),
    .X(clknet_1_0__leaf_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net281 (.A(clknet_0_net281),
    .X(clknet_1_1__leaf_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net280 (.A(net280),
    .X(clknet_0_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net280 (.A(clknet_0_net280),
    .X(clknet_1_0__leaf_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net280 (.A(clknet_0_net280),
    .X(clknet_1_1__leaf_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net654 (.A(net654),
    .X(clknet_0_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net654 (.A(clknet_0_net654),
    .X(clknet_1_0__leaf_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net654 (.A(clknet_0_net654),
    .X(clknet_1_1__leaf_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net855 (.A(net855),
    .X(clknet_0_net855));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net855 (.A(clknet_0_net855),
    .X(clknet_1_0__leaf_net855));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net855 (.A(clknet_0_net855),
    .X(clknet_1_1__leaf_net855));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net404 (.A(net404),
    .X(clknet_0_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net404 (.A(clknet_0_net404),
    .X(clknet_1_0__leaf_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net404 (.A(clknet_0_net404),
    .X(clknet_1_1__leaf_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net859 (.A(net859),
    .X(clknet_0_net859));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net859 (.A(clknet_0_net859),
    .X(clknet_1_0__leaf_net859));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net859 (.A(clknet_0_net859),
    .X(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net874 (.A(net874),
    .X(clknet_0_net874));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net874 (.A(clknet_0_net874),
    .X(clknet_1_0__leaf_net874));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net874 (.A(clknet_0_net874),
    .X(clknet_1_1__leaf_net874));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net196 (.A(net196),
    .X(clknet_0_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net196 (.A(clknet_0_net196),
    .X(clknet_1_0__leaf_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net196 (.A(clknet_0_net196),
    .X(clknet_1_1__leaf_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net156 (.A(net156),
    .X(clknet_0_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net156 (.A(clknet_0_net156),
    .X(clknet_1_0__leaf_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net156 (.A(clknet_0_net156),
    .X(clknet_1_1__leaf_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net155 (.A(net155),
    .X(clknet_0_net155));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net155 (.A(clknet_0_net155),
    .X(clknet_1_0__leaf_net155));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net155 (.A(clknet_0_net155),
    .X(clknet_1_1__leaf_net155));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net130 (.A(net130),
    .X(clknet_0_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net130 (.A(clknet_0_net130),
    .X(clknet_1_0__leaf_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net130 (.A(clknet_0_net130),
    .X(clknet_1_1__leaf_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net375 (.A(net375),
    .X(clknet_0_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net375 (.A(clknet_0_net375),
    .X(clknet_1_0__leaf_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net375 (.A(clknet_0_net375),
    .X(clknet_1_1__leaf_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net373 (.A(net373),
    .X(clknet_0_net373));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net373 (.A(clknet_0_net373),
    .X(clknet_1_0__leaf_net373));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net373 (.A(clknet_0_net373),
    .X(clknet_1_1__leaf_net373));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net217),
    .X(net910));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer2 (.A(net910),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net1003),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net217),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net86),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net914),
    .X(net915));
 sky130_fd_sc_hd__buf_4 rebuffer7 (.A(net675),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net916),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net917),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net85),
    .X(net919));
 sky130_fd_sc_hd__clkbuf_2 rebuffer11 (.A(net423),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net920),
    .X(net921));
 sky130_fd_sc_hd__clkbuf_1 rebuffer13 (.A(net921),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net70),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net421),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net438),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net925),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net438),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net438),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net211),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net436),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net930),
    .X(net931));
 sky130_fd_sc_hd__buf_2 rebuffer23 (.A(net436),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net932),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net932),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net934),
    .X(net935));
 sky130_fd_sc_hd__buf_6 rebuffer27 (.A(net421),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(net424),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net204),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(net938),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer31 (.A(net203),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(net203),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(net941),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net678),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net339),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net803),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net260),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net699),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net42),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net55),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net469),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net322),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net124),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net679),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net171),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net166),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net323),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net349),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net685),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net344),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net707),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net568),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net565),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net363),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net303),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net123),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net708),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net325),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net495),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net498),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net509),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net324),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net192),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net750),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net321),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net400),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net713),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net429),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net447),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net596),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net669),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net458),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net854),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net297),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net693),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net696),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net715),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net387),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net710),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net419),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net744),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net271),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net667),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net650),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net877),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net714),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net143),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net479),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net670),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(net685),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net316),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net714),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(net684),
    .X(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_X (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_D (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_B1_N (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_RESET_B (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_B (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_D (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_X (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_SCD (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_X (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A3 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A3 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_X (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_B1_N (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_Q_N (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A0 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_Q (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A3 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_D (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_SCE (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_X (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_Y (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A0 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_RESET_B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_SET_B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A3 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_S1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_X (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_SCD (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_B1_N (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_X (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_SET_B (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_X (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_D (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_SCE (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_SCD (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_X (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_X (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_RESET_B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A0 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A4 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_SCE (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_Y (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_Y (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_B1_N (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_S1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_S0 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B1_N (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_Y (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_X (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_B1_N (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A0 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A3 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_SCE (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_X (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_S0 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_B (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A3 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_SCE (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_Q (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer4_A (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer3_A (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_A (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_RESET_B (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_RESET_B (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_D (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_X (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A3 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_Y (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_S0 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_D (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_B1_N (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_SCE (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_D (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_SCE (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_D (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_SCE (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A3 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_B1_N (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_Y (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A0 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_S0 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_SCD (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_D (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_Q (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A0 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S0 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_RESET_B (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_SCE (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S0 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_RESET_B (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_RESET_B (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_X (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A3 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_RESET_B (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_X (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_SCD (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A3 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_S0 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_SCE (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_RESET_B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_X (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A2 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_SCD (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_SET_B (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A4 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A3 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_Q (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_B1_N (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_SCE (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_S1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_Q_N (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_Q (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_D (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_SET_B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_SCD (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A3 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_SCD (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_SCD (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_X (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S0 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A0 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_SET_B (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A3 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_X (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_A3 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_X (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_RESET_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S0 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A0 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A0 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_X (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_A3 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_Y (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A0 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A3 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S0 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_SCE (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A3 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S0 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_B (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_X (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A0 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_SCE (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_X (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_Y (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap124_A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A3 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A4 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_D (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_B (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_Y (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_S0 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_D (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_SET_B (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_SCE (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_D (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_SCD (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_SCE (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_X (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A3 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_B1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_S1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_SET_B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S0 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_RESET_B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_Y (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A3 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c653_A1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c652_A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_A1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_S0 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_B (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_B (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_Q (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c640_A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_SET_B (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A0 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_B (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_Y (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_SET_B (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_D (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_SCD (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_SET_B (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A3 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A3 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_SCD (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_SCD (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_Y (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold35_A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_SCE (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_A3 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_Q (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A0 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_S1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_S0 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A3 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A2 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_X (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_B1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_RESET_B (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A0 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A3 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A3 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_Y (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_D (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_RESET_B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A2 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A4 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_Y (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_B1_N (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_Q_N (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_RESET_B (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_D (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A3 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_Q (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A3 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A1 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S0 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S1 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_B1 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_X (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_D (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A1 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_X (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A0 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A3 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_RESET_B (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A1 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A3 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A1 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_B1 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_X (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_RESET_B (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_SCE (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_B1_N (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A0 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_Q (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_D (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_X (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_D (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_SCD (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_B (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_S1 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_Y (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_X (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap120_A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c657_DE (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_D (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_S0 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_Y (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_D (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_D (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_SET_B (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_X (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A0 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_SCE (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_RESET_B (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_SCD (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_X (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_SCD (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_Q_N (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A0 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_Q (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_B1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A3 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_Q_N (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A0 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_B1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A3 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A3 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_Q (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_D (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_S1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_SCD (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_X (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge740_S0 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A0 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A2 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_D (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_Y (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A2 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A1 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A2 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A0 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_RESET_B (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_SET_B (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_X (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S0 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A0 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A2 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_SCE (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A2 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A2 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_X (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_D (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A2 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_SCD (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A2 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_S1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_X (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A0 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_X (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A2 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A2 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_SCD (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_X (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A3 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_SCD (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c652_B1_N (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c648_A3 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_S0 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c641_A (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c638_Y (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A0 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_S0 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A0 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_SCD (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c657_SCD (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_SCE (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c640_Y (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A3 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A3 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c648_A2 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_A1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_SCD (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c645_B (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_A2 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c643_Q (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A2 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_S1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_D (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_S0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_RESET_B (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c649_S1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_X (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A0 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A3 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_SCE (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_B1 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_X (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A0 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A1 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A1 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_X (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A2 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_S1 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_s745_Q (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net672_A (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_s763_GCLK (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold44_A (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_s772_Q (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S0 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A4 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A3 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c650_S0 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A3 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A3 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_S1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B1_N (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B1_N (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_Y (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_s787_Q (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S0 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_SET_B (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_B1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_X (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_D (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A3 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_S0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_SET_B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B1_N (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_X (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_s835_Q (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S0 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S0 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S0 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_SCD (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A4 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_SCD (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_X (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A3 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A3 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_Y (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_SCD (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_B1_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A3 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A3 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A3 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_RESET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_X (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A2 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A1 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A2 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_RESET_B (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A2 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_B1_N (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A2 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_B1_N (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A3 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_B (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_B (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_B1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_B (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A3 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A2 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S0 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A2 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A0 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_B1_N (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_S1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_B (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S0 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_B1_N (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A2 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_B1_N (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A2 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A2 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_A1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_SCD (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_A2 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_D (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_RESET_B (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_A3 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A4 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A3 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A2 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S0 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A1 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_A1 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A2 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_S1 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_B1 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A0 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A4 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A0 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A3 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B1_N (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_B1_N (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_B (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_SCE (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A3 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B1 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_B (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_SCE (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A2 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A2 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A2 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A3 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A2 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_S0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_S0 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_B (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_B1_N (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A2 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A3 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_SCE (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_B1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_A2 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_A3 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A2 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A0 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_B1_N (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_SET_B (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SCE (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold36_A (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_A3 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_X (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A0 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_SCE (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_A0 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_SCE (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A3 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_B1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_D (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_X (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A0 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A2 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A2 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A3 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A3 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_X (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_B1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A3 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A3 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B1_N (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A3 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_SET_B (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A2 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_X (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_SCD (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A3 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A2 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_SET_B (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A2 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_SET_B (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_X (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_SCD (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_SET_B (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A3 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_X (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_B (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A3 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_B (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_RESET_B (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_SET_B (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_X (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_SET_B (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_SCD (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A3 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_A3 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_B (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_Q (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A3 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A2 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_X (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_Q (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_X (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_Q (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A3 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_X (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A1 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A3 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A1 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A3 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_B1_N (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_X (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A3 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A2 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A2 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_X (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A2 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_Q (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_X (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net859_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_s746_GCLK (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_s742_Q (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_S1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_s752_Q (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A3 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_B1 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_B1_N (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_X (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A3 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A3 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A3 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_S0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A2 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_SET_B (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_SCE (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_S0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap120_X (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A1 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A0 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_S1 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A3 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_X (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A3 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_D (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A3 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_S0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_SCD (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_X (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A0 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_DE (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A4 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_S0 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c658_SCE (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_SCD (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c653_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_DE (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A2 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_X (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_X (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A0 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A3 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A3 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A3 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S0 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A3 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A3 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_S0 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_B1_N (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A0 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_X (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_B (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A2 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B1_N (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A4 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_B1_N (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_B1_N (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_B1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_S1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B1_N (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_X (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A0 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A3 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S0 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A0 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A3 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A3 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_X (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_D (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A3 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_RESET_B (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A2 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_SET_B (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A4 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap129_X (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_SCE (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_RESET_B (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A2 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_RESET_B (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_RESET_B (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_SCD (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_B (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap131_X (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_D (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_A2 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_B1_N (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_B1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_X (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_RESET_B (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A4 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_A3 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_DE (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_A4 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_B (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_X (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_SCE (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_B1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_SCE (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_SET_B (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_SET_B (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_S1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A3 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_X (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_S1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_S1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_SCE (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_SCE (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_SET_B (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A3 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_X (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_S0 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_SCD (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A2 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_SCE (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A2 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A3 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A2 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A2 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap137_X (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_D (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B1_N (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_RESET_B (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_B (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_S0 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_X (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_RESET_B (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A4 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_SET_B (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B1_N (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_B (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_A2 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_A3 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_SCE (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A4 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A2 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_B1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_SCD (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_SCD (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_SET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_S1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_X (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S0 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_X (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_B1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S0 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_SET_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_SET_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_B1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B1_N (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S0 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_S1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_S1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_X (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_SCD (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_A4 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_B1_N (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_A2 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_A2 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A3 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_B (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_B (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_X (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A4 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A4 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A4 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A3 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_X (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_SCD (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_SCE (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A3 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_B1_N (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_X (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S0 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S0 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_SCE (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A3 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_B1_N (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A3 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A2 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_X (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_B1_N (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_B1_N (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A2 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B1_N (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_S0 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_X (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_RESET_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_S0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_SCD (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_D (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_SCE (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_X (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_S0 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A1 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A2 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A2 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A2 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_B1_N (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_CLK_N (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_X (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_X (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_X (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_X (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_B1 (.DIODE(clknet_1_0__leaf_net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_B1 (.DIODE(clknet_1_0__leaf_net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_S1 (.DIODE(clknet_1_0__leaf_net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S0 (.DIODE(clknet_1_0__leaf_net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_S0 (.DIODE(clknet_1_0__leaf_net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net716_X (.DIODE(clknet_1_0__leaf_net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A2 (.DIODE(clknet_1_0__leaf_net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_RESET_B (.DIODE(clknet_1_0__leaf_net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A3 (.DIODE(clknet_1_0__leaf_net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net576_X (.DIODE(clknet_1_0__leaf_net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S1 (.DIODE(clknet_1_1__leaf_net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(clknet_1_1__leaf_net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net834_X (.DIODE(clknet_1_1__leaf_net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S0 (.DIODE(clknet_1_0__leaf_net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_SCE (.DIODE(clknet_1_0__leaf_net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_SCE (.DIODE(clknet_1_0__leaf_net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A3 (.DIODE(clknet_1_0__leaf_net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A3 (.DIODE(clknet_1_0__leaf_net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net826_X (.DIODE(clknet_1_0__leaf_net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_SCD (.DIODE(clknet_1_1__leaf_net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(clknet_1_1__leaf_net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net826_X (.DIODE(clknet_1_1__leaf_net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_SCE (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_B1 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_RESET_B (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A2 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A3 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A3 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_B1_N (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A3 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A4 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A3 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A3 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net386_X (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_S1 (.DIODE(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A0 (.DIODE(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S0 (.DIODE(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A2 (.DIODE(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A0 (.DIODE(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S0 (.DIODE(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A0 (.DIODE(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net386_X (.DIODE(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_S1 (.DIODE(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_S0 (.DIODE(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_S1 (.DIODE(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S1 (.DIODE(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_B1_N (.DIODE(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net655_X (.DIODE(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S1 (.DIODE(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_SET_B (.DIODE(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S1 (.DIODE(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_SCD (.DIODE(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A3 (.DIODE(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S0 (.DIODE(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net655_X (.DIODE(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(clknet_1_1__leaf_net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(clknet_1_1__leaf_net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net855_X (.DIODE(clknet_1_1__leaf_net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S1 (.DIODE(clknet_1_0__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_S0 (.DIODE(clknet_1_0__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_B1_N (.DIODE(clknet_1_0__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_SET_B (.DIODE(clknet_1_0__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_S1 (.DIODE(clknet_1_0__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net859_X (.DIODE(clknet_1_0__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_B1 (.DIODE(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_S1 (.DIODE(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_SCE (.DIODE(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S0 (.DIODE(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A4 (.DIODE(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net859_X (.DIODE(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_SCE (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_X (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer14_X (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer20_X (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer25_A (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer24_A (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_SCD (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A2 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer23_X (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net873));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(net217),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer35 (.A(net1003),
    .X(net1004));
 sky130_fd_sc_hd__mux4_1 clone36 (.A0(net216),
    .A1(net215),
    .A2(net213),
    .A3(net201),
    .S0(net896),
    .S1(net207),
    .X(net1005));
 sky130_fd_sc_hd__clkbuf_1 clone37 (.A(net1007),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer38 (.A(net199),
    .X(net1007));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
