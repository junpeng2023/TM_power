module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in3,
    in4,
    in5,
    in6,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out3,
    out4,
    out5,
    out6,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in3;
 input in4;
 input in5;
 input in6;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out3;
 output out4;
 output out5;
 output out6;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_0_net527;
 wire clknet_1_0__leaf_net527;
 wire clknet_1_1__leaf_net527;
 wire clknet_0_net627;
 wire clknet_1_0__leaf_net627;
 wire clknet_1_1__leaf_net627;
 wire clknet_0_net652;
 wire clknet_1_0__leaf_net652;
 wire clknet_1_1__leaf_net652;
 wire clknet_0_net629;
 wire clknet_1_0__leaf_net629;
 wire clknet_1_1__leaf_net629;
 wire clknet_0_net620;
 wire clknet_1_0__leaf_net620;
 wire clknet_1_1__leaf_net620;
 wire clknet_0_net656;
 wire clknet_1_0__leaf_net656;
 wire clknet_1_1__leaf_net656;
 wire clknet_0_net524;
 wire clknet_1_0__leaf_net524;
 wire clknet_1_1__leaf_net524;
 wire clknet_0_net517;
 wire clknet_1_0__leaf_net517;
 wire clknet_1_1__leaf_net517;
 wire clknet_0_net523;
 wire clknet_1_0__leaf_net523;
 wire clknet_1_1__leaf_net523;
 wire clknet_0_net525;
 wire clknet_1_0__leaf_net525;
 wire clknet_1_1__leaf_net525;
 wire clknet_0_net519;
 wire clknet_1_0__leaf_net519;
 wire clknet_1_1__leaf_net519;
 wire clknet_0_net569;
 wire clknet_1_0__leaf_net569;
 wire clknet_1_1__leaf_net569;
 wire clknet_0_net508;
 wire clknet_1_0__leaf_net508;
 wire clknet_1_1__leaf_net508;
 wire clknet_0_net511;
 wire clknet_1_0__leaf_net511;
 wire clknet_1_1__leaf_net511;
 wire clknet_0_net396;
 wire clknet_1_0__leaf_net396;
 wire clknet_1_1__leaf_net396;
 wire clknet_0_net518;
 wire clknet_1_0__leaf_net518;
 wire clknet_1_1__leaf_net518;
 wire clknet_0_net398;
 wire clknet_1_0__leaf_net398;
 wire clknet_1_1__leaf_net398;
 wire clknet_0_net337;
 wire clknet_1_0__leaf_net337;
 wire clknet_1_1__leaf_net337;
 wire clknet_0_net465;
 wire clknet_1_0__leaf_net465;
 wire clknet_1_1__leaf_net465;
 wire clknet_0_net800;
 wire clknet_1_0__leaf_net800;
 wire clknet_1_1__leaf_net800;
 wire clknet_0_net452;
 wire clknet_1_0__leaf_net452;
 wire clknet_1_1__leaf_net452;
 wire clknet_0_net333;
 wire clknet_1_0__leaf_net333;
 wire clknet_1_1__leaf_net333;
 wire clknet_0_net797;
 wire clknet_1_0__leaf_net797;
 wire clknet_1_1__leaf_net797;
 wire clknet_0_net229;
 wire clknet_1_0__leaf_net229;
 wire clknet_1_1__leaf_net229;
 wire clknet_0_net221;
 wire clknet_1_0__leaf_net221;
 wire clknet_1_1__leaf_net221;
 wire clknet_0_net142;
 wire clknet_1_0__leaf_net142;
 wire clknet_1_1__leaf_net142;
 wire clknet_0_net423;
 wire clknet_1_0__leaf_net423;
 wire clknet_1_1__leaf_net423;
 wire clknet_0_net575;
 wire clknet_1_0__leaf_net575;
 wire clknet_1_1__leaf_net575;
 wire clknet_0_net272;
 wire clknet_1_0__leaf_net272;
 wire clknet_1_1__leaf_net272;
 wire clknet_0_net150;
 wire clknet_1_0__leaf_net150;
 wire clknet_1_1__leaf_net150;
 wire clknet_0_net140;
 wire clknet_1_0__leaf_net140;
 wire clknet_1_1__leaf_net140;
 wire clknet_0_net149;
 wire clknet_1_0__leaf_net149;
 wire clknet_1_1__leaf_net149;
 wire clknet_0_net301;
 wire clknet_1_0__leaf_net301;
 wire clknet_1_1__leaf_net301;
 wire clknet_0_net429;
 wire clknet_1_0__leaf_net429;
 wire clknet_1_1__leaf_net429;
 wire clknet_0_net308;
 wire clknet_1_0__leaf_net308;
 wire clknet_1_1__leaf_net308;
 wire clknet_0_net300;
 wire clknet_1_0__leaf_net300;
 wire clknet_1_1__leaf_net300;
 wire clknet_0_net595;
 wire clknet_1_0__leaf_net595;
 wire clknet_1_1__leaf_net595;
 wire clknet_0_net449;
 wire clknet_1_0__leaf_net449;
 wire clknet_1_1__leaf_net449;
 wire clknet_0_net153;
 wire clknet_1_0__leaf_net153;
 wire clknet_1_1__leaf_net153;
 wire clknet_0_net151;
 wire clknet_1_0__leaf_net151;
 wire clknet_1_1__leaf_net151;
 wire clknet_0_net306;
 wire clknet_1_0__leaf_net306;
 wire clknet_1_1__leaf_net306;
 wire clknet_0_net298;
 wire clknet_1_0__leaf_net298;
 wire clknet_1_1__leaf_net298;
 wire clknet_0_net784;
 wire clknet_1_0__leaf_net784;
 wire clknet_1_1__leaf_net784;
 wire clknet_0_net135;
 wire clknet_1_0__leaf_net135;
 wire clknet_1_1__leaf_net135;
 wire clknet_0_net277;
 wire clknet_1_0__leaf_net277;
 wire clknet_1_1__leaf_net277;
 wire clknet_0_net334;
 wire clknet_1_0__leaf_net334;
 wire clknet_1_1__leaf_net334;
 wire clknet_0_net336;
 wire clknet_1_0__leaf_net336;
 wire clknet_1_1__leaf_net336;
 wire clknet_0_net335;
 wire clknet_1_0__leaf_net335;
 wire clknet_1_1__leaf_net335;
 wire clknet_0_net287;
 wire clknet_1_0__leaf_net287;
 wire clknet_1_1__leaf_net287;
 wire clknet_0_net405;
 wire clknet_1_0__leaf_net405;
 wire clknet_1_1__leaf_net405;
 wire clknet_0_net290;
 wire clknet_1_0__leaf_net290;
 wire clknet_1_1__leaf_net290;
 wire clknet_0_net129;
 wire clknet_1_0__leaf_net129;
 wire clknet_1_1__leaf_net129;
 wire clknet_0_net621;
 wire clknet_1_0__leaf_net621;
 wire clknet_1_1__leaf_net621;
 wire clknet_0_net130;
 wire clknet_1_0__leaf_net130;
 wire clknet_1_1__leaf_net130;
 wire clknet_0_net387;
 wire clknet_1_0__leaf_net387;
 wire clknet_1_1__leaf_net387;
 wire clknet_0_net393;
 wire clknet_1_0__leaf_net393;
 wire clknet_1_1__leaf_net393;
 wire clknet_0_net789;
 wire clknet_1_0__leaf_net789;
 wire clknet_1_1__leaf_net789;
 wire clknet_0_net162;
 wire clknet_1_0__leaf_net162;
 wire clknet_1_1__leaf_net162;
 wire clknet_0_net156;
 wire clknet_1_0__leaf_net156;
 wire clknet_1_1__leaf_net156;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;

 sky130_fd_sc_hd__and2_0 c100 (.A(net70),
    .B(net85),
    .X(net87));
 sky130_fd_sc_hd__and2_0 c101 (.A(net86),
    .B(net87),
    .X(net88));
 sky130_fd_sc_hd__mux4_1 c102 (.A0(net10),
    .A1(net88),
    .A2(net86),
    .A3(net83),
    .S0(net70),
    .S1(net38),
    .X(net89));
 sky130_fd_sc_hd__dlrtn_1 c103 (.D(net76),
    .GATE_N(clknet_leaf_9_clk),
    .RESET_B(net78),
    .Q(net90));
 sky130_fd_sc_hd__and3_1 c104 (.A(net9),
    .B(net85),
    .C(net83),
    .X(net91));
 sky130_fd_sc_hd__dlrtn_1 c105 (.D(net49),
    .GATE_N(clknet_leaf_8_clk),
    .RESET_B(net76),
    .Q(net92));
 sky130_fd_sc_hd__and2_1 c106 (.A(net75),
    .B(net3),
    .X(net93));
 sky130_fd_sc_hd__dlrtp_1 c107 (.D(net76),
    .GATE(clknet_leaf_8_clk),
    .RESET_B(net52),
    .Q(net94));
 sky130_fd_sc_hd__dlrtp_1 c108 (.D(net15),
    .GATE(clknet_leaf_8_clk),
    .RESET_B(net93),
    .Q(net95));
 sky130_fd_sc_hd__dlrtp_1 c109 (.D(net829),
    .GATE(clknet_leaf_9_clk),
    .RESET_B(net57),
    .Q(net96));
 sky130_fd_sc_hd__and2_0 c110 (.A(net873),
    .B(net83),
    .X(net97));
 sky130_fd_sc_hd__mux4_1 c111 (.A0(net94),
    .A1(net40),
    .A2(net93),
    .A3(net75),
    .S0(net37),
    .S1(net26),
    .X(net98));
 sky130_fd_sc_hd__edfxbp_1 c112 (.CLK(clknet_leaf_9_clk),
    .D(net93),
    .DE(net887),
    .Q(net791),
    .Q_N(net99));
 sky130_fd_sc_hd__and2_1 c113 (.A(net95),
    .B(net75),
    .X(net100));
 sky130_fd_sc_hd__and2_0 c114 (.A(net79),
    .B(net40),
    .X(net101));
 sky130_fd_sc_hd__and2_0 c115 (.A(net79),
    .B(net732),
    .X(net102));
 sky130_fd_sc_hd__and2_0 c116 (.A(net52),
    .B(net760),
    .X(net103));
 sky130_fd_sc_hd__and2_0 c117 (.A(net103),
    .B(net101),
    .X(net104));
 sky130_fd_sc_hd__and3_1 c118 (.A(net83),
    .B(net95),
    .C(net100),
    .X(net105));
 sky130_fd_sc_hd__dfbbn_1 c119 (.CLK_N(clknet_leaf_8_clk),
    .D(net105),
    .RESET_B(net95),
    .SET_B(net93),
    .Q(net107),
    .Q_N(net106));
 sky130_fd_sc_hd__and2_0 c120 (.A(net107),
    .B(net101),
    .X(net108));
 sky130_fd_sc_hd__dfbbp_1 c121 (.CLK(clknet_leaf_8_clk),
    .D(net102),
    .RESET_B(net108),
    .SET_B(net106),
    .Q(net110),
    .Q_N(net109));
 sky130_fd_sc_hd__edfxtp_1 c122 (.CLK(clknet_leaf_8_clk),
    .D(net108),
    .DE(net93),
    .Q(net782));
 sky130_fd_sc_hd__and2_0 c123 (.A(net92),
    .B(net109),
    .X(net111));
 sky130_fd_sc_hd__sdfxbp_1 c124 (.CLK(clknet_leaf_8_clk),
    .D(net904),
    .SCD(net107),
    .SCE(net105),
    .Q(net112));
 sky130_fd_sc_hd__and2_1 c125 (.A(net111),
    .B(net112),
    .X(net113));
 sky130_fd_sc_hd__buf_1 c126 (.A(net772),
    .X(net114));
 sky130_fd_sc_hd__buf_1 c127 (.A(net114),
    .X(net115));
 sky130_fd_sc_hd__and2_1 c128 (.A(net764),
    .B(net758),
    .X(net116));
 sky130_fd_sc_hd__buf_1 c129 (.A(net757),
    .X(net117));
 sky130_fd_sc_hd__buf_1 c130 (.A(net117),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 c131 (.A(net776),
    .X(net119));
 sky130_fd_sc_hd__and2_2 c132 (.A(net759),
    .B(net117),
    .X(net120));
 sky130_fd_sc_hd__and2_2 c133 (.A(net119),
    .B(net758),
    .X(net121));
 sky130_fd_sc_hd__and2_1 c134 (.A(net773),
    .B(net803),
    .X(net122));
 sky130_fd_sc_hd__and2_2 c135 (.A(net116),
    .B(net120),
    .X(net123));
 sky130_fd_sc_hd__and2_2 c136 (.A(net122),
    .B(net119),
    .X(net124));
 sky130_fd_sc_hd__dfxtp_2 c137 (.CLK(clknet_leaf_0_clk),
    .D(net123),
    .Q(net125));
 sky130_fd_sc_hd__and2_2 c138 (.A(net759),
    .B(net118),
    .X(net126));
 sky130_fd_sc_hd__and2_4 c139 (.A(net767),
    .B(net754),
    .X(net127));
 sky130_fd_sc_hd__buf_2 c140 (.A(net124),
    .X(net128));
 sky130_fd_sc_hd__sdlclkp_1 c141 (.CLK(clknet_leaf_26_clk),
    .GATE(net118),
    .SCE(net128),
    .GCLK(net129));
 sky130_fd_sc_hd__and2_0 c142 (.A(net125),
    .B(clknet_1_1__leaf_net129),
    .X(net130));
 sky130_fd_sc_hd__mux4_1 c143 (.A0(net128),
    .A1(net116),
    .A2(net772),
    .A3(net754),
    .S0(net114),
    .S1(net124),
    .X(net131));
 sky130_fd_sc_hd__and2_4 c144 (.A(net115),
    .B(net834),
    .X(net132));
 sky130_fd_sc_hd__sdfxbp_1 c145 (.CLK(clknet_leaf_6_clk),
    .D(net754),
    .SCD(clknet_1_0__leaf_net130),
    .SCE(net132),
    .Q(net134),
    .Q_N(net133));
 sky130_fd_sc_hd__sdlclkp_2 c146 (.CLK(clknet_leaf_4_clk),
    .GATE(net870),
    .SCE(net132),
    .GCLK(net135));
 sky130_fd_sc_hd__and2_0 c147 (.A(net127),
    .B(net6),
    .X(net136));
 sky130_fd_sc_hd__buf_1 c148 (.A(net136),
    .X(net137));
 sky130_fd_sc_hd__buf_1 c149 (.A(net0),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_2 c150 (.A(net114),
    .X(net139));
 sky130_fd_sc_hd__dlclkp_1 c151 (.CLK(clknet_leaf_0_clk),
    .GATE(net123),
    .GCLK(net140));
 sky130_fd_sc_hd__buf_2 c152 (.A(net770),
    .X(net141));
 sky130_fd_sc_hd__sdlclkp_4 c153 (.CLK(clknet_leaf_5_clk),
    .GATE(net137),
    .SCE(net0),
    .GCLK(net142));
 sky130_fd_sc_hd__buf_2 c154 (.A(net120),
    .X(net143));
 sky130_fd_sc_hd__and2_2 c155 (.A(net762),
    .B(net121),
    .X(net144));
 sky130_fd_sc_hd__and2_0 c156 (.A(net139),
    .B(clknet_1_1__leaf_net140),
    .X(net784));
 sky130_fd_sc_hd__dlymetal6s2s_1 c157 (.A(net141),
    .X(net145));
 sky130_fd_sc_hd__and2_1 c158 (.A(net758),
    .B(net11),
    .X(net146));
 sky130_fd_sc_hd__and2_2 c159 (.A(net138),
    .B(net803),
    .X(net147));
 sky130_fd_sc_hd__and2_1 c160 (.A(net136),
    .B(net6),
    .X(net148));
 sky130_fd_sc_hd__buf_1 c161 (.A(clknet_1_0__leaf_net140),
    .X(net149));
 sky130_fd_sc_hd__and2_0 c162 (.A(clknet_1_1__leaf_net142),
    .B(net120),
    .X(net150));
 sky130_fd_sc_hd__buf_1 c163 (.A(clknet_1_0__leaf_net149),
    .X(net151));
 sky130_fd_sc_hd__sdfxtp_2 c164 (.CLK(clknet_leaf_5_clk),
    .D(clknet_1_0__leaf_net151),
    .SCD(net137),
    .SCE(net769),
    .Q(net152));
 sky130_fd_sc_hd__and3_1 c165 (.A(net152),
    .B(clknet_1_1__leaf_net151),
    .C(clknet_1_1__leaf_net149),
    .X(net153));
 sky130_fd_sc_hd__dfrbp_1 c166 (.CLK(clknet_leaf_1_clk),
    .D(net148),
    .RESET_B(net816),
    .Q(net155),
    .Q_N(net154));
 sky130_fd_sc_hd__and3_1 c167 (.A(net6),
    .B(clknet_1_0__leaf_net130),
    .C(net154),
    .X(net156));
 sky130_fd_sc_hd__and2_0 c168 (.A(net778),
    .B(clknet_1_0__leaf_net130),
    .X(net789));
 sky130_fd_sc_hd__and2_4 c169 (.A(net41),
    .B(net866),
    .X(net157));
 sky130_fd_sc_hd__dfrbp_1 c170 (.CLK(clknet_leaf_14_clk),
    .D(net754),
    .RESET_B(net144),
    .Q(net159),
    .Q_N(net158));
 sky130_fd_sc_hd__sdfxtp_2 c171 (.CLK(clknet_leaf_1_clk),
    .D(clknet_1_0__leaf_net140),
    .SCD(net148),
    .SCE(net28),
    .Q(net160));
 sky130_fd_sc_hd__and2_1 c172 (.A(net825),
    .B(net124),
    .X(net161));
 sky130_fd_sc_hd__and3_1 c173 (.A(clknet_1_0__leaf_net789),
    .B(net116),
    .C(net803),
    .X(net162));
 sky130_fd_sc_hd__dfrtn_1 c174 (.CLK_N(clknet_leaf_6_clk),
    .D(net756),
    .RESET_B(net157),
    .Q(net163));
 sky130_fd_sc_hd__and2_0 c175 (.A(net146),
    .B(net121),
    .X(net164));
 sky130_fd_sc_hd__dfrtp_1 c176 (.CLK(clknet_leaf_12_clk),
    .D(net144),
    .RESET_B(clknet_1_1__leaf_net162),
    .Q(net165));
 sky130_fd_sc_hd__dfrtp_4 c177 (.CLK(clknet_leaf_0_clk),
    .D(net126),
    .RESET_B(net817),
    .Q(net166));
 sky130_fd_sc_hd__dfrtp_1 c178 (.CLK(clknet_leaf_5_clk),
    .D(net148),
    .RESET_B(net24),
    .Q(net167));
 sky130_fd_sc_hd__and3_2 c179 (.A(net0),
    .B(net33),
    .C(net29),
    .X(net168));
 sky130_fd_sc_hd__dfsbp_1 c180 (.CLK(clknet_leaf_14_clk),
    .D(net23),
    .SET_B(net12),
    .Q(net170),
    .Q_N(net169));
 sky130_fd_sc_hd__and2_1 c181 (.A(net757),
    .B(net809),
    .X(net171));
 sky130_fd_sc_hd__dfsbp_1 c182 (.CLK(clknet_leaf_12_clk),
    .D(net171),
    .SET_B(net161),
    .Q(net173),
    .Q_N(net172));
 sky130_fd_sc_hd__and2_1 c183 (.A(net159),
    .B(net169),
    .X(net174));
 sky130_fd_sc_hd__dfstp_1 c184 (.CLK(clknet_leaf_12_clk),
    .D(net857),
    .SET_B(net157),
    .Q(net175));
 sky130_fd_sc_hd__and2_0 c185 (.A(net760),
    .B(net166),
    .X(net176));
 sky130_fd_sc_hd__dfstp_1 c186 (.CLK(clknet_leaf_18_clk),
    .D(net164),
    .SET_B(net141),
    .Q(net177));
 sky130_fd_sc_hd__and3_1 c187 (.A(net174),
    .B(net172),
    .C(net7),
    .X(net178));
 sky130_fd_sc_hd__dfstp_1 c188 (.CLK(clknet_leaf_5_clk),
    .D(net137),
    .SET_B(net821),
    .Q(net179));
 sky130_fd_sc_hd__and2_1 c189 (.A(net60),
    .B(net768),
    .X(net180));
 sky130_fd_sc_hd__and2_1 c190 (.A(net773),
    .B(net761),
    .X(net181));
 sky130_fd_sc_hd__and2_1 c191 (.A(net774),
    .B(net733),
    .X(net182));
 sky130_fd_sc_hd__dlrbn_1 c192 (.D(net870),
    .GATE_N(clknet_leaf_12_clk),
    .RESET_B(clknet_1_0__leaf_net153),
    .Q(net184),
    .Q_N(net183));
 sky130_fd_sc_hd__and2_0 c193 (.A(net159),
    .B(net183),
    .X(net185));
 sky130_fd_sc_hd__and2_0 c194 (.A(net167),
    .B(net28),
    .X(net186));
 sky130_fd_sc_hd__dlrbn_1 c195 (.D(net164),
    .GATE_N(clknet_leaf_18_clk),
    .RESET_B(net143),
    .Q(net188),
    .Q_N(net187));
 sky130_fd_sc_hd__and2_1 c196 (.A(net122),
    .B(net180),
    .X(net189));
 sky130_fd_sc_hd__and2_1 c197 (.A(net61),
    .B(net183),
    .X(net190));
 sky130_fd_sc_hd__dlrbp_1 c198 (.D(net161),
    .GATE(clknet_leaf_4_clk),
    .RESET_B(net38),
    .Q(net192),
    .Q_N(net191));
 sky130_fd_sc_hd__and2_2 c199 (.A(net20),
    .B(net189),
    .X(net790));
 sky130_fd_sc_hd__and2_0 c200 (.A(net775),
    .B(net61),
    .X(net193));
 sky130_fd_sc_hd__and2_2 c201 (.A(net185),
    .B(net767),
    .X(net194));
 sky130_fd_sc_hd__and2_1 c202 (.A(net181),
    .B(net191),
    .X(net195));
 sky130_fd_sc_hd__and2_1 c203 (.A(net192),
    .B(net195),
    .X(net196));
 sky130_fd_sc_hd__and2_1 c204 (.A(net189),
    .B(net158),
    .X(net197));
 sky130_fd_sc_hd__and2_0 c205 (.A(net193),
    .B(net174),
    .X(net198));
 sky130_fd_sc_hd__and2_2 c206 (.A(net188),
    .B(net11),
    .X(net802));
 sky130_fd_sc_hd__dlrbp_1 c207 (.D(net198),
    .GATE(clknet_leaf_14_clk),
    .RESET_B(net802),
    .Q(net200),
    .Q_N(net199));
 sky130_fd_sc_hd__and2_0 c208 (.A(net843),
    .B(net177),
    .X(net201));
 sky130_fd_sc_hd__and2_1 c209 (.A(net844),
    .B(net193),
    .X(net202));
 sky130_fd_sc_hd__and2_1 c210 (.A(net78),
    .B(net194),
    .X(net203));
 sky130_fd_sc_hd__dlrtn_1 c211 (.D(net809),
    .GATE_N(clknet_leaf_14_clk),
    .RESET_B(net202),
    .Q(net204));
 sky130_fd_sc_hd__dlrtn_1 c212 (.D(net178),
    .GATE_N(clknet_leaf_10_clk),
    .RESET_B(net817),
    .Q(net205));
 sky130_fd_sc_hd__and2_0 c213 (.A(net38),
    .B(net26),
    .X(net206));
 sky130_fd_sc_hd__dlrtn_1 c214 (.D(net88),
    .GATE_N(clknet_leaf_10_clk),
    .RESET_B(net802),
    .Q(net207));
 sky130_fd_sc_hd__sdfrbp_1 c215 (.CLK(clknet_leaf_6_clk),
    .D(net882),
    .RESET_B(net202),
    .SCD(net770),
    .SCE(net803),
    .Q(net209),
    .Q_N(net208));
 sky130_fd_sc_hd__and2_0 c216 (.A(net205),
    .B(net766),
    .X(net210));
 sky130_fd_sc_hd__dlrtp_1 c217 (.D(net73),
    .GATE(clknet_leaf_10_clk),
    .RESET_B(clknet_1_0__leaf_net784),
    .Q(net211));
 sky130_fd_sc_hd__dlrtp_1 c218 (.D(net174),
    .GATE(clknet_leaf_7_clk),
    .RESET_B(net57),
    .Q(net212));
 sky130_fd_sc_hd__dlrtp_1 c219 (.D(net186),
    .GATE(clknet_leaf_5_clk),
    .RESET_B(net82),
    .Q(net213));
 sky130_fd_sc_hd__and2_1 c220 (.A(net87),
    .B(net865),
    .X(net214));
 sky130_fd_sc_hd__edfxbp_1 c221 (.CLK(clknet_leaf_12_clk),
    .D(net29),
    .DE(net178),
    .Q(net215));
 sky130_fd_sc_hd__sdfxtp_1 c222 (.CLK(clknet_leaf_7_clk),
    .D(net202),
    .SCD(net895),
    .SCE(net29),
    .Q(net216));
 sky130_fd_sc_hd__and2_1 c223 (.A(net213),
    .B(net208),
    .X(net217));
 sky130_fd_sc_hd__edfxtp_1 c224 (.CLK(clknet_leaf_20_clk),
    .D(net82),
    .DE(net147),
    .Q(net218));
 sky130_fd_sc_hd__and2_1 c225 (.A(net209),
    .B(net160),
    .X(net219));
 sky130_fd_sc_hd__and2_0 c226 (.A(net66),
    .B(net8),
    .X(net220));
 sky130_fd_sc_hd__sdlclkp_1 c227 (.CLK(clknet_leaf_7_clk),
    .GATE(net846),
    .SCE(net57),
    .GCLK(net221));
 sky130_fd_sc_hd__and2_1 c228 (.A(net27),
    .B(net218),
    .X(net222));
 sky130_fd_sc_hd__and2_0 c229 (.A(net865),
    .B(net220),
    .X(net223));
 sky130_fd_sc_hd__or4bb_1 c230 (.A(net212),
    .B(net216),
    .C_N(clknet_1_0__leaf_net221),
    .D_N(net127),
    .X(net224));
 sky130_fd_sc_hd__and2_0 c231 (.A(net113),
    .B(net774),
    .X(net225));
 sky130_fd_sc_hd__and2_0 c232 (.A(net875),
    .B(net113),
    .X(net226));
 sky130_fd_sc_hd__dfbbn_1 c233 (.CLK_N(clknet_leaf_10_clk),
    .D(net42),
    .RESET_B(net145),
    .SET_B(net100),
    .Q(net227));
 sky130_fd_sc_hd__and2_0 c234 (.A(net227),
    .B(net206),
    .X(net228));
 sky130_fd_sc_hd__dfbbn_1 c235 (.CLK_N(clknet_leaf_9_clk),
    .D(net104),
    .RESET_B(net67),
    .SET_B(net754),
    .Q(net781));
 sky130_fd_sc_hd__sdlclkp_2 c236 (.CLK(clknet_leaf_9_clk),
    .GATE(net57),
    .SCE(net104),
    .GCLK(net229));
 sky130_fd_sc_hd__and2_1 c237 (.A(net817),
    .B(net37),
    .X(net230));
 sky130_fd_sc_hd__dfbbp_1 c238 (.CLK(clknet_leaf_10_clk),
    .D(net64),
    .RESET_B(net207),
    .SET_B(net194),
    .Q(net231));
 sky130_fd_sc_hd__sdfxbp_1 c239 (.CLK(clknet_leaf_15_clk),
    .D(net100),
    .SCD(clknet_1_1__leaf_net153),
    .SCE(net230),
    .Q(net232));
 sky130_fd_sc_hd__and3_1 c240 (.A(net232),
    .B(net204),
    .C(clknet_1_0__leaf_net229),
    .X(net233));
 sky130_fd_sc_hd__and2_0 c241 (.A(net754),
    .B(net16),
    .X(net234));
 sky130_fd_sc_hd__and3_1 c242 (.A(net190),
    .B(net771),
    .C(net230),
    .X(net235));
 sky130_fd_sc_hd__and2_0 c243 (.A(net204),
    .B(net2),
    .X(net236));
 sky130_fd_sc_hd__and2_0 c244 (.A(net206),
    .B(net84),
    .X(net237));
 sky130_fd_sc_hd__sdlclkp_4 c245 (.CLK(clknet_leaf_16_clk),
    .GATE(net236),
    .SCE(net210),
    .GCLK(net797));
 sky130_fd_sc_hd__sdfxbp_1 c246 (.CLK(clknet_leaf_11_clk),
    .D(net225),
    .SCD(net207),
    .SCE(net790),
    .Q(net239),
    .Q_N(net238));
 sky130_fd_sc_hd__sdfxtp_1 c247 (.CLK(clknet_leaf_9_clk),
    .D(net97),
    .SCD(net908),
    .SCE(net100),
    .Q(net240));
 sky130_fd_sc_hd__and3_1 c248 (.A(net180),
    .B(net190),
    .C(clknet_1_0__leaf_net229),
    .X(net241));
 sky130_fd_sc_hd__sdfxtp_1 c249 (.CLK(clknet_leaf_10_clk),
    .D(net3),
    .SCD(net113),
    .SCE(net64),
    .Q(net242));
 sky130_fd_sc_hd__clkbuf_2 c25 (.A(net770),
    .X(net0));
 sky130_fd_sc_hd__dfrbp_1 c250 (.CLK(clknet_leaf_11_clk),
    .D(net234),
    .RESET_B(net235),
    .Q(net243));
 sky130_fd_sc_hd__dfrbp_1 c251 (.CLK(clknet_leaf_11_clk),
    .D(net241),
    .RESET_B(net814),
    .Q(net245),
    .Q_N(net244));
 sky130_fd_sc_hd__clkbuf_4 c252 (.A(net121),
    .X(net246));
 sky130_fd_sc_hd__dfrtn_1 c253 (.CLK_N(clknet_leaf_0_clk),
    .D(net126),
    .RESET_B(net246),
    .Q(net247));
 sky130_fd_sc_hd__buf_1 c254 (.A(net778),
    .X(net248));
 sky130_fd_sc_hd__and2_1 c255 (.A(net762),
    .B(net118),
    .X(net249));
 sky130_fd_sc_hd__and2_1 c256 (.A(net247),
    .B(net755),
    .X(net250));
 sky130_fd_sc_hd__and2_2 c257 (.A(net250),
    .B(net122),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 c258 (.A(net122),
    .X(net252));
 sky130_fd_sc_hd__dfrtp_2 c259 (.CLK(clknet_leaf_25_clk),
    .D(net251),
    .RESET_B(net128),
    .Q(net253));
 sky130_fd_sc_hd__clkbuf_4 c26 (.A(net775),
    .X(net1));
 sky130_fd_sc_hd__dfrtp_1 c260 (.CLK(clknet_leaf_33_clk),
    .D(net755),
    .RESET_B(net246),
    .Q(net254));
 sky130_fd_sc_hd__buf_1 c261 (.A(net765),
    .X(net255));
 sky130_fd_sc_hd__dfrtp_2 c262 (.CLK(clknet_leaf_1_clk),
    .D(net255),
    .RESET_B(net132),
    .Q(net256));
 sky130_fd_sc_hd__and2_1 c263 (.A(net114),
    .B(net248),
    .X(net257));
 sky130_fd_sc_hd__and2_1 c264 (.A(net253),
    .B(net247),
    .X(net258));
 sky130_fd_sc_hd__sdfxtp_1 c265 (.CLK(clknet_leaf_32_clk),
    .D(net763),
    .SCD(net890),
    .SCE(net246),
    .Q(net259));
 sky130_fd_sc_hd__clkbuf_1 c266 (.A(net254),
    .X(net260));
 sky130_fd_sc_hd__and2_1 c267 (.A(net876),
    .B(net250),
    .X(net261));
 sky130_fd_sc_hd__and3_1 c268 (.A(net260),
    .B(net256),
    .C(net762),
    .X(net262));
 sky130_fd_sc_hd__and2_2 c269 (.A(net257),
    .B(net260),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_2 c27 (.A(net1),
    .X(net2));
 sky130_fd_sc_hd__dfsbp_1 c270 (.CLK(clknet_leaf_30_clk),
    .D(net263),
    .SET_B(net261),
    .Q(net265),
    .Q_N(net264));
 sky130_fd_sc_hd__dfsbp_2 c271 (.CLK(clknet_leaf_29_clk),
    .D(net261),
    .SET_B(net263),
    .Q(net267),
    .Q_N(net266));
 sky130_fd_sc_hd__and3_1 c272 (.A(net248),
    .B(net258),
    .C(net849),
    .X(net268));
 sky130_fd_sc_hd__dfstp_1 c273 (.CLK(clknet_leaf_0_clk),
    .D(net246),
    .SET_B(net123),
    .Q(net269));
 sky130_fd_sc_hd__and2_1 c274 (.A(net5),
    .B(net255),
    .X(net270));
 sky130_fd_sc_hd__dfstp_2 c275 (.CLK(clknet_leaf_24_clk),
    .D(net147),
    .SET_B(net773),
    .Q(net271));
 sky130_fd_sc_hd__and3_1 c276 (.A(net252),
    .B(clknet_1_1__leaf_net142),
    .C(net146),
    .X(net272));
 sky130_fd_sc_hd__and2_1 c277 (.A(net146),
    .B(net757),
    .X(net273));
 sky130_fd_sc_hd__dfstp_4 c278 (.CLK(clknet_leaf_5_clk),
    .D(net767),
    .SET_B(clknet_1_0__leaf_net272),
    .Q(net274));
 sky130_fd_sc_hd__dfbbn_1 c279 (.CLK_N(clknet_leaf_13_clk),
    .D(net758),
    .RESET_B(net273),
    .SET_B(net146),
    .Q(net276),
    .Q_N(net275));
 sky130_fd_sc_hd__clkbuf_2 c28 (.A(net8),
    .X(net3));
 sky130_fd_sc_hd__and2_0 c280 (.A(clknet_1_0__leaf_net135),
    .B(net17),
    .X(net277));
 sky130_fd_sc_hd__and2_0 c281 (.A(net772),
    .B(net17),
    .X(net278));
 sky130_fd_sc_hd__and2_1 c282 (.A(net764),
    .B(net4),
    .X(net279));
 sky130_fd_sc_hd__dlrbn_1 c283 (.D(net252),
    .GATE_N(clknet_leaf_13_clk),
    .RESET_B(net263),
    .Q(net281),
    .Q_N(net280));
 sky130_fd_sc_hd__and2_2 c284 (.A(net278),
    .B(net270),
    .X(net282));
 sky130_fd_sc_hd__dlrbn_1 c285 (.D(net260),
    .GATE_N(clknet_leaf_29_clk),
    .RESET_B(net282),
    .Q(net284),
    .Q_N(net283));
 sky130_fd_sc_hd__dfbbn_1 c286 (.CLK_N(clknet_leaf_21_clk),
    .D(net270),
    .RESET_B(net144),
    .SET_B(net840),
    .Q(net286),
    .Q_N(net285));
 sky130_fd_sc_hd__and2_0 c287 (.A(net284),
    .B(clknet_1_0__leaf_net277),
    .X(net287));
 sky130_fd_sc_hd__dlrbp_1 c288 (.D(net282),
    .GATE(clknet_leaf_13_clk),
    .RESET_B(net271),
    .Q(net289),
    .Q_N(net288));
 sky130_fd_sc_hd__and2_0 c289 (.A(clknet_1_1__leaf_net287),
    .B(net757),
    .X(net290));
 sky130_fd_sc_hd__and2_1 c29 (.A(net1),
    .B(net0),
    .X(net4));
 sky130_fd_sc_hd__dlrbp_1 c290 (.D(net273),
    .GATE(clknet_leaf_4_clk),
    .RESET_B(net279),
    .Q(net292),
    .Q_N(net291));
 sky130_fd_sc_hd__and2_2 c291 (.A(net289),
    .B(net280),
    .X(net783));
 sky130_fd_sc_hd__dlrtn_1 c292 (.D(net862),
    .GATE_N(clknet_leaf_4_clk),
    .RESET_B(net246),
    .Q(net293));
 sky130_fd_sc_hd__dfbbp_1 c293 (.CLK(clknet_leaf_13_clk),
    .D(clknet_1_1__leaf_net272),
    .RESET_B(net855),
    .SET_B(net282),
    .Q(net295),
    .Q_N(net294));
 sky130_fd_sc_hd__dlrtn_1 c294 (.D(net279),
    .GATE_N(clknet_leaf_6_clk),
    .RESET_B(net163),
    .Q(net296));
 sky130_fd_sc_hd__and2_0 c295 (.A(net296),
    .B(net155),
    .X(net297));
 sky130_fd_sc_hd__and2_0 c296 (.A(clknet_1_1__leaf_net151),
    .B(net774),
    .X(net298));
 sky130_fd_sc_hd__and2_0 c297 (.A(net278),
    .B(net285),
    .X(net299));
 sky130_fd_sc_hd__and2_0 c298 (.A(clknet_1_1__leaf_net149),
    .B(net274),
    .X(net300));
 sky130_fd_sc_hd__and2_0 c299 (.A(net163),
    .B(clknet_1_1__leaf_net149),
    .X(net301));
 sky130_fd_sc_hd__and2_1 c30 (.A(net771),
    .B(net763),
    .X(net5));
 sky130_fd_sc_hd__sdfxbp_1 c300 (.CLK(clknet_leaf_4_clk),
    .D(net273),
    .SCD(net293),
    .SCE(clknet_1_1__leaf_net300),
    .Q(net303),
    .Q_N(net302));
 sky130_fd_sc_hd__dlrtn_1 c301 (.D(net857),
    .GATE_N(clknet_leaf_12_clk),
    .RESET_B(net157),
    .Q(net304));
 sky130_fd_sc_hd__dlrtp_1 c302 (.D(net176),
    .GATE(clknet_leaf_12_clk),
    .RESET_B(clknet_1_0__leaf_net162),
    .Q(net305));
 sky130_fd_sc_hd__and2_0 c303 (.A(net4),
    .B(clknet_1_0__leaf_net151),
    .X(net306));
 sky130_fd_sc_hd__and2_0 c304 (.A(net119),
    .B(net771),
    .X(net307));
 sky130_fd_sc_hd__a2111o_1 c305 (.A1(clknet_1_1__leaf_net301),
    .A2(net291),
    .B1(net778),
    .C1(net33),
    .D1(net305),
    .X(net308));
 sky130_fd_sc_hd__mux4_1 c306 (.A0(net179),
    .A1(net296),
    .A2(net33),
    .A3(clknet_1_0__leaf_net149),
    .S0(clknet_1_0__leaf_net308),
    .S1(net758),
    .X(net309));
 sky130_fd_sc_hd__dlrtp_1 c307 (.D(clknet_1_0__leaf_net272),
    .GATE(clknet_leaf_4_clk),
    .RESET_B(clknet_1_1__leaf_net306),
    .Q(net310));
 sky130_fd_sc_hd__dlrtp_2 c308 (.D(clknet_1_0__leaf_net306),
    .GATE(clknet_leaf_5_clk),
    .RESET_B(clknet_1_0__leaf_net150),
    .Q(net311));
 sky130_fd_sc_hd__a2111o_1 c309 (.A1(net171),
    .A2(net31),
    .B1(net310),
    .C1(net116),
    .D1(net302),
    .X(net312));
 sky130_fd_sc_hd__buf_1 c31 (.A(net754),
    .X(net6));
 sky130_fd_sc_hd__and2_0 c310 (.A(net296),
    .B(net311),
    .X(net313));
 sky130_fd_sc_hd__edfxbp_1 c311 (.CLK(clknet_leaf_6_clk),
    .D(net313),
    .DE(clknet_1_1__leaf_net308),
    .Q(net314));
 sky130_fd_sc_hd__edfxtp_1 c312 (.CLK(clknet_leaf_4_clk),
    .D(net33),
    .DE(net22),
    .Q(net315));
 sky130_fd_sc_hd__sdfxbp_1 c313 (.CLK(clknet_leaf_5_clk),
    .D(net297),
    .SCD(net893),
    .SCE(net157),
    .Q(net317),
    .Q_N(net316));
 sky130_fd_sc_hd__and2_2 c314 (.A(net313),
    .B(net316),
    .X(net318));
 sky130_fd_sc_hd__and2_0 c315 (.A(net281),
    .B(net51),
    .X(net319));
 sky130_fd_sc_hd__and2_2 c316 (.A(net318),
    .B(net319),
    .X(net320));
 sky130_fd_sc_hd__sdfxtp_2 c317 (.CLK(clknet_leaf_14_clk),
    .D(net11),
    .SCD(net145),
    .SCE(net197),
    .Q(net321));
 sky130_fd_sc_hd__mux4_1 c318 (.A0(net320),
    .A1(net24),
    .A2(net768),
    .A3(net321),
    .S0(net311),
    .S1(net274),
    .X(net322));
 sky130_fd_sc_hd__or4bb_4 c319 (.A(net317),
    .B(net267),
    .C_N(net900),
    .D_N(net11),
    .X(net323));
 sky130_fd_sc_hd__and2_2 c32 (.A(net770),
    .B(net5),
    .X(net7));
 sky130_fd_sc_hd__sdfxtp_1 c320 (.CLK(clknet_leaf_14_clk),
    .D(net825),
    .SCD(clknet_1_1__leaf_net290),
    .SCE(net189),
    .Q(net324));
 sky130_fd_sc_hd__and2_0 c321 (.A(net319),
    .B(net39),
    .X(net325));
 sky130_fd_sc_hd__mux4_1 c322 (.A0(net307),
    .A1(clknet_1_0__leaf_net290),
    .A2(net775),
    .A3(net275),
    .S0(net182),
    .S1(net194),
    .X(net326));
 sky130_fd_sc_hd__sdlclkp_1 c323 (.CLK(clknet_leaf_14_clk),
    .GATE(net293),
    .SCE(net157),
    .GCLK(net327));
 sky130_fd_sc_hd__and3_1 c324 (.A(net44),
    .B(net321),
    .C(net315),
    .X(net328));
 sky130_fd_sc_hd__and2_1 c325 (.A(net303),
    .B(net163),
    .X(net329));
 sky130_fd_sc_hd__and2_1 c326 (.A(net305),
    .B(net35),
    .X(net330));
 sky130_fd_sc_hd__sdlclkp_2 c327 (.CLK(clknet_leaf_14_clk),
    .GATE(net328),
    .SCE(clknet_1_1__leaf_net300),
    .GCLK(net800));
 sky130_fd_sc_hd__sdfbbn_1 c328 (.CLK_N(clknet_leaf_17_clk),
    .D(clknet_1_0__leaf_net800),
    .RESET_B(net320),
    .SCD(net323),
    .SCE(net194),
    .SET_B(net839),
    .Q(net332),
    .Q_N(net331));
 sky130_fd_sc_hd__and3_1 c329 (.A(net329),
    .B(clknet_1_0__leaf_net800),
    .C(net293),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_4 c33 (.A(net756),
    .X(net8));
 sky130_fd_sc_hd__and2_0 c330 (.A(clknet_1_1__leaf_net277),
    .B(net737),
    .X(net334));
 sky130_fd_sc_hd__and2_0 c331 (.A(clknet_1_0__leaf_net334),
    .B(net44),
    .X(net335));
 sky130_fd_sc_hd__and2_0 c332 (.A(net321),
    .B(clknet_1_1__leaf_net334),
    .X(net336));
 sky130_fd_sc_hd__sdlclkp_4 c333 (.CLK(clknet_leaf_17_clk),
    .GATE(clknet_1_1__leaf_net336),
    .SCE(net331),
    .GCLK(net337));
 sky130_fd_sc_hd__and2_0 c334 (.A(net286),
    .B(net125),
    .X(net338));
 sky130_fd_sc_hd__dfrbp_2 c335 (.CLK(clknet_leaf_17_clk),
    .D(net338),
    .RESET_B(clknet_1_0__leaf_net336),
    .Q(net799),
    .Q_N(net339));
 sky130_fd_sc_hd__and2_0 c336 (.A(net759),
    .B(net731),
    .X(net340));
 sky130_fd_sc_hd__mux4_1 c337 (.A0(clknet_1_0__leaf_net162),
    .A1(net269),
    .A2(net251),
    .A3(net21),
    .S0(net764),
    .S1(net736),
    .X(net341));
 sky130_fd_sc_hd__sdfrtn_1 c338 (.CLK_N(clknet_leaf_15_clk),
    .D(net165),
    .RESET_B(net22),
    .SCD(net802),
    .SCE(clknet_1_1__leaf_net300),
    .Q(net342));
 sky130_fd_sc_hd__and3_1 c339 (.A(net735),
    .B(net166),
    .C(net267),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_2 c34 (.A(net5),
    .X(net9));
 sky130_fd_sc_hd__and3_1 c340 (.A(net276),
    .B(net175),
    .C(clknet_1_0__leaf_net789),
    .X(net344));
 sky130_fd_sc_hd__sdfxtp_1 c341 (.CLK(clknet_leaf_14_clk),
    .D(net344),
    .SCD(net219),
    .SCE(net342),
    .Q(net345));
 sky130_fd_sc_hd__and3_1 c342 (.A(net894),
    .B(net340),
    .C(net736),
    .X(net346));
 sky130_fd_sc_hd__and2_0 c343 (.A(net218),
    .B(net56),
    .X(net347));
 sky130_fd_sc_hd__and3_1 c344 (.A(net345),
    .B(net276),
    .C(net343),
    .X(net348));
 sky130_fd_sc_hd__dfbbn_1 c345 (.CLK_N(clknet_leaf_17_clk),
    .D(net197),
    .RESET_B(net139),
    .SET_B(net315),
    .Q(net350),
    .Q_N(net349));
 sky130_fd_sc_hd__and2_0 c346 (.A(net71),
    .B(net820),
    .X(net351));
 sky130_fd_sc_hd__and3_1 c347 (.A(net175),
    .B(net325),
    .C(net71),
    .X(net352));
 sky130_fd_sc_hd__and2_0 c348 (.A(net70),
    .B(net735),
    .X(net353));
 sky130_fd_sc_hd__dfbbn_1 c349 (.CLK_N(clknet_leaf_12_clk),
    .D(net883),
    .RESET_B(net352),
    .SET_B(net832),
    .Q(net355),
    .Q_N(net354));
 sky130_fd_sc_hd__and2_2 c35 (.A(net6),
    .B(net9),
    .X(net10));
 sky130_fd_sc_hd__and3_1 c350 (.A(net332),
    .B(net349),
    .C(net730),
    .X(net356));
 sky130_fd_sc_hd__sdfbbp_1 c351 (.CLK(clknet_leaf_12_clk),
    .D(net69),
    .RESET_B(clknet_1_1__leaf_net162),
    .SCD(net354),
    .SCE(net896),
    .SET_B(net808),
    .Q(net357));
 sky130_fd_sc_hd__and3_4 c352 (.A(net343),
    .B(net80),
    .C(net310),
    .X(net358));
 sky130_fd_sc_hd__and3_1 c353 (.A(net81),
    .B(net802),
    .C(net353),
    .X(net359));
 sky130_fd_sc_hd__and3_1 c354 (.A(net763),
    .B(net358),
    .C(net269),
    .X(net360));
 sky130_fd_sc_hd__dfbbp_1 c355 (.CLK(clknet_leaf_11_clk),
    .D(net223),
    .RESET_B(net320),
    .SET_B(net358),
    .Q(net361));
 sky130_fd_sc_hd__and3_1 c356 (.A(net342),
    .B(net361),
    .C(net85),
    .X(net362));
 sky130_fd_sc_hd__and2_0 c357 (.A(net330),
    .B(clknet_1_0__leaf_net135),
    .X(net363));
 sky130_fd_sc_hd__and3_1 c358 (.A(net84),
    .B(net245),
    .C(net766),
    .X(net801));
 sky130_fd_sc_hd__dfrbp_1 c359 (.CLK(clknet_leaf_16_clk),
    .D(net766),
    .RESET_B(clknet_1_1__leaf_net153),
    .Q(net365),
    .Q_N(net364));
 sky130_fd_sc_hd__and2_1 c36 (.A(net758),
    .B(net760),
    .X(net11));
 sky130_fd_sc_hd__and3_1 c360 (.A(net355),
    .B(net86),
    .C(net238),
    .X(net795));
 sky130_fd_sc_hd__and3_1 c361 (.A(clknet_1_1__leaf_net129),
    .B(clknet_1_1__leaf_net221),
    .C(net365),
    .X(net366));
 sky130_fd_sc_hd__sdfxbp_1 c362 (.CLK(clknet_leaf_16_clk),
    .D(net210),
    .SCD(net68),
    .SCE(net350),
    .Q(net367));
 sky130_fd_sc_hd__and2_0 c363 (.A(net876),
    .B(net145),
    .X(net368));
 sky130_fd_sc_hd__sdfxbp_1 c364 (.CLK(clknet_leaf_10_clk),
    .D(net836),
    .SCD(net359),
    .SCE(net330),
    .Q(net369));
 sky130_fd_sc_hd__and2_1 c365 (.A(net771),
    .B(net340),
    .X(net779));
 sky130_fd_sc_hd__a2111o_1 c366 (.A1(net230),
    .A2(net369),
    .B1(net86),
    .C1(net364),
    .D1(net760),
    .X(net370));
 sky130_fd_sc_hd__and2_0 c367 (.A(net56),
    .B(net350),
    .X(net371));
 sky130_fd_sc_hd__sdfrtp_1 c368 (.CLK(clknet_leaf_10_clk),
    .D(clknet_1_1__leaf_net135),
    .RESET_B(net808),
    .SCD(clknet_1_0__leaf_net335),
    .SCE(clknet_1_1__leaf_net129),
    .Q(net372));
 sky130_fd_sc_hd__and2_0 c369 (.A(net327),
    .B(net219),
    .X(net373));
 sky130_fd_sc_hd__and2_4 c37 (.A(net772),
    .B(net2),
    .X(net12));
 sky130_fd_sc_hd__and3_1 c370 (.A(net370),
    .B(net373),
    .C(net244),
    .X(net374));
 sky130_fd_sc_hd__and2_0 c371 (.A(net184),
    .B(net237),
    .X(net375));
 sky130_fd_sc_hd__and2_0 c372 (.A(net372),
    .B(net231),
    .X(net786));
 sky130_fd_sc_hd__sdfxtp_1 c373 (.CLK(clknet_leaf_15_clk),
    .D(net374),
    .SCD(net362),
    .SCE(net783),
    .Q(net376));
 sky130_fd_sc_hd__dfrtn_1 c374 (.CLK_N(clknet_leaf_16_clk),
    .D(net367),
    .RESET_B(clknet_1_1__leaf_net335),
    .Q(net377));
 sky130_fd_sc_hd__dfrtp_1 c375 (.CLK(clknet_leaf_15_clk),
    .D(net368),
    .RESET_B(net351),
    .Q(net378));
 sky130_fd_sc_hd__and3_1 c376 (.A(net377),
    .B(net378),
    .C(net85),
    .X(net787));
 sky130_fd_sc_hd__and3_1 c377 (.A(net228),
    .B(net233),
    .C(net787),
    .X(net379));
 sky130_fd_sc_hd__and2_1 c378 (.A(net776),
    .B(net766),
    .X(net380));
 sky130_fd_sc_hd__buf_1 c379 (.A(net380),
    .X(net381));
 sky130_fd_sc_hd__and2_2 c38 (.A(net11),
    .B(net771),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 c380 (.A(net776),
    .X(net382));
 sky130_fd_sc_hd__and2_1 c381 (.A(net259),
    .B(net254),
    .X(net383));
 sky130_fd_sc_hd__dlymetal6s2s_1 c382 (.A(net382),
    .X(net384));
 sky130_fd_sc_hd__buf_1 c383 (.A(net760),
    .X(net385));
 sky130_fd_sc_hd__dlymetal6s2s_1 c384 (.A(net759),
    .X(net386));
 sky130_fd_sc_hd__and2_0 c385 (.A(net763),
    .B(clknet_1_1__leaf_net130),
    .X(net387));
 sky130_fd_sc_hd__dlymetal6s2s_1 c386 (.A(net383),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_2 c387 (.A(net772),
    .X(net389));
 sky130_fd_sc_hd__sdfxtp_1 c388 (.CLK(clknet_leaf_27_clk),
    .D(net384),
    .SCD(net251),
    .SCE(net263),
    .Q(net390));
 sky130_fd_sc_hd__clkbuf_1 c389 (.A(net385),
    .X(net391));
 sky130_fd_sc_hd__dfrbp_1 c39 (.CLK(clknet_leaf_7_clk),
    .D(net2),
    .RESET_B(net12),
    .Q(net15),
    .Q_N(net14));
 sky130_fd_sc_hd__and2_1 c390 (.A(net247),
    .B(net388),
    .X(net392));
 sky130_fd_sc_hd__and2_0 c391 (.A(net391),
    .B(clknet_1_1__leaf_net387),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_2 c392 (.A(net268),
    .X(net394));
 sky130_fd_sc_hd__dfrtp_1 c393 (.CLK(clknet_leaf_27_clk),
    .D(net392),
    .RESET_B(net384),
    .Q(net395));
 sky130_fd_sc_hd__dlclkp_2 c394 (.CLK(clknet_leaf_26_clk),
    .GATE(clknet_1_0__leaf_net393),
    .GCLK(net396));
 sky130_fd_sc_hd__dfrtp_4 c395 (.CLK(clknet_leaf_33_clk),
    .D(net123),
    .RESET_B(net831),
    .Q(net397));
 sky130_fd_sc_hd__and3_1 c396 (.A(net395),
    .B(clknet_1_1__leaf_net396),
    .C(clknet_1_0__leaf_net387),
    .X(net398));
 sky130_fd_sc_hd__sdfxtp_1 c397 (.CLK(clknet_leaf_32_clk),
    .D(clknet_1_0__leaf_net398),
    .SCD(net383),
    .SCE(net901),
    .Q(net399));
 sky130_fd_sc_hd__and3_2 c398 (.A(net397),
    .B(net390),
    .C(net399),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_2 c399 (.A(net729),
    .X(net401));
 sky130_fd_sc_hd__and2_4 c40 (.A(net903),
    .B(net8),
    .X(net16));
 sky130_fd_sc_hd__buf_1 c400 (.A(net891),
    .X(net402));
 sky130_fd_sc_hd__dfsbp_1 c401 (.CLK(clknet_leaf_3_clk),
    .D(net5),
    .SET_B(net394),
    .Q(net404),
    .Q_N(net403));
 sky130_fd_sc_hd__and2_0 c402 (.A(clknet_1_0__leaf_net287),
    .B(clknet_1_1__leaf_net156),
    .X(net405));
 sky130_fd_sc_hd__and2_1 c403 (.A(net269),
    .B(net1),
    .X(net406));
 sky130_fd_sc_hd__dfsbp_1 c404 (.CLK(clknet_leaf_27_clk),
    .D(net392),
    .SET_B(net282),
    .Q(net408),
    .Q_N(net407));
 sky130_fd_sc_hd__and3_1 c405 (.A(net382),
    .B(net261),
    .C(net837),
    .X(net409));
 sky130_fd_sc_hd__and2_1 c406 (.A(net127),
    .B(net402),
    .X(net410));
 sky130_fd_sc_hd__dfstp_1 c407 (.CLK(clknet_leaf_32_clk),
    .D(net263),
    .SET_B(net822),
    .Q(net411));
 sky130_fd_sc_hd__and2_1 c408 (.A(net406),
    .B(net774),
    .X(net412));
 sky130_fd_sc_hd__and2_1 c409 (.A(net391),
    .B(net138),
    .X(net413));
 sky130_fd_sc_hd__dfxbp_1 c41 (.CLK(clknet_leaf_3_clk),
    .D(net12),
    .Q(net18),
    .Q_N(net17));
 sky130_fd_sc_hd__dfbbn_1 c410 (.CLK_N(clknet_leaf_29_clk),
    .D(net413),
    .RESET_B(net115),
    .SET_B(net294),
    .Q(net415),
    .Q_N(net414));
 sky130_fd_sc_hd__and2_1 c411 (.A(net253),
    .B(net400),
    .X(net416));
 sky130_fd_sc_hd__dfstp_1 c412 (.CLK(clknet_leaf_22_clk),
    .D(net402),
    .SET_B(net123),
    .Q(net417));
 sky130_fd_sc_hd__dfstp_1 c413 (.CLK(clknet_leaf_24_clk),
    .D(net410),
    .SET_B(net413),
    .Q(net418));
 sky130_fd_sc_hd__dlrbn_1 c414 (.D(clknet_1_1__leaf_net405),
    .GATE_N(clknet_leaf_22_clk),
    .RESET_B(clknet_1_0__leaf_net387),
    .Q(net420),
    .Q_N(net419));
 sky130_fd_sc_hd__dlrbn_1 c415 (.D(net282),
    .GATE_N(clknet_leaf_29_clk),
    .RESET_B(clknet_1_0__leaf_net156),
    .Q(net422),
    .Q_N(net421));
 sky130_fd_sc_hd__and2_0 c416 (.A(net418),
    .B(clknet_1_0__leaf_net142),
    .X(net423));
 sky130_fd_sc_hd__dfbbn_1 c417 (.CLK_N(clknet_leaf_24_clk),
    .D(net417),
    .RESET_B(net147),
    .SET_B(net410),
    .Q(net425),
    .Q_N(net424));
 sky130_fd_sc_hd__dfbbp_1 c418 (.CLK(clknet_leaf_0_clk),
    .D(net837),
    .RESET_B(net807),
    .SET_B(clknet_1_0__leaf_net398),
    .Q(net427),
    .Q_N(net426));
 sky130_fd_sc_hd__and3_1 c419 (.A(net420),
    .B(net417),
    .C(net424),
    .X(net428));
 sky130_fd_sc_hd__dfxbp_1 c42 (.CLK(clknet_leaf_7_clk),
    .D(net10),
    .Q(net20),
    .Q_N(net19));
 sky130_fd_sc_hd__and3_1 c420 (.A(net769),
    .B(net17),
    .C(clknet_1_1__leaf_net301),
    .X(net429));
 sky130_fd_sc_hd__mux4_1 c421 (.A0(net765),
    .A1(net37),
    .A2(net139),
    .A3(clknet_1_1__leaf_net429),
    .S0(net380),
    .S1(net803),
    .X(net430));
 sky130_fd_sc_hd__sdfxbp_1 c422 (.CLK(clknet_leaf_3_clk),
    .D(net116),
    .SCD(clknet_1_0__leaf_net429),
    .SCE(net22),
    .Q(net432),
    .Q_N(net431));
 sky130_fd_sc_hd__and2_0 c423 (.A(net755),
    .B(net312),
    .X(net433));
 sky130_fd_sc_hd__dlrbp_1 c424 (.D(net433),
    .GATE(clknet_leaf_3_clk),
    .RESET_B(net431),
    .Q(net434));
 sky130_fd_sc_hd__and2_0 c425 (.A(net170),
    .B(net769),
    .X(net435));
 sky130_fd_sc_hd__and2_0 c426 (.A(net289),
    .B(net21),
    .X(net436));
 sky130_fd_sc_hd__and2_2 c427 (.A(net18),
    .B(net758),
    .X(net796));
 sky130_fd_sc_hd__and2_0 c428 (.A(net312),
    .B(net761),
    .X(net437));
 sky130_fd_sc_hd__and2_1 c429 (.A(net436),
    .B(net7),
    .X(net438));
 sky130_fd_sc_hd__buf_1 c43 (.A(net803),
    .X(net21));
 sky130_fd_sc_hd__and2_1 c430 (.A(net297),
    .B(net154),
    .X(net439));
 sky130_fd_sc_hd__dlrbp_1 c431 (.D(clknet_1_0__leaf_net306),
    .GATE(clknet_leaf_1_clk),
    .RESET_B(net879),
    .Q(net441),
    .Q_N(net440));
 sky130_fd_sc_hd__sdfxbp_1 c432 (.CLK(clknet_leaf_21_clk),
    .D(net438),
    .SCD(net796),
    .SCE(net421),
    .Q(net443),
    .Q_N(net442));
 sky130_fd_sc_hd__sdfxtp_1 c433 (.CLK(clknet_leaf_3_clk),
    .D(net437),
    .SCD(net863),
    .SCE(net120),
    .Q(net444));
 sky130_fd_sc_hd__and2_2 c434 (.A(net441),
    .B(net269),
    .X(net445));
 sky130_fd_sc_hd__and3_1 c435 (.A(net434),
    .B(net436),
    .C(net444),
    .X(net446));
 sky130_fd_sc_hd__and3_1 c436 (.A(net155),
    .B(net442),
    .C(net445),
    .X(net447));
 sky130_fd_sc_hd__and2_1 c437 (.A(net443),
    .B(net447),
    .X(net448));
 sky130_fd_sc_hd__and3_1 c438 (.A(net383),
    .B(clknet_1_0__leaf_net300),
    .C(net31),
    .X(net449));
 sky130_fd_sc_hd__dlrtn_1 c439 (.D(net435),
    .GATE_N(clknet_leaf_26_clk),
    .RESET_B(clknet_1_0__leaf_net449),
    .Q(net450));
 sky130_fd_sc_hd__and2_2 c44 (.A(net758),
    .B(net3),
    .X(net22));
 sky130_fd_sc_hd__sdfxtp_1 c440 (.CLK(clknet_leaf_26_clk),
    .D(clknet_1_0__leaf_net449),
    .SCD(net251),
    .SCE(net450),
    .Q(net451));
 sky130_fd_sc_hd__and3_1 c441 (.A(net23),
    .B(net796),
    .C(clknet_1_0__leaf_net800),
    .X(net452));
 sky130_fd_sc_hd__and3_1 c442 (.A(net54),
    .B(net323),
    .C(net739),
    .X(net453));
 sky130_fd_sc_hd__sdfxtp_1 c443 (.CLK(clknet_leaf_18_clk),
    .D(clknet_1_1__leaf_net130),
    .SCD(clknet_1_1__leaf_net452),
    .SCE(net453),
    .Q(net454));
 sky130_fd_sc_hd__or4bb_2 c444 (.A(net53),
    .B(net295),
    .C_N(net189),
    .D_N(net274),
    .X(net455));
 sky130_fd_sc_hd__and2_1 c445 (.A(net415),
    .B(net262),
    .X(net456));
 sky130_fd_sc_hd__sdfbbn_1 c446 (.CLK_N(clknet_leaf_18_clk),
    .D(net324),
    .RESET_B(net810),
    .SCD(net790),
    .SCE(net315),
    .SET_B(clknet_1_1__leaf_net452),
    .Q(net457));
 sky130_fd_sc_hd__dfbbn_1 c447 (.CLK_N(clknet_leaf_13_clk),
    .D(clknet_1_0__leaf_net290),
    .RESET_B(clknet_1_0__leaf_net452),
    .SET_B(net53),
    .Q(net459),
    .Q_N(net458));
 sky130_fd_sc_hd__dfbbn_1 c448 (.CLK_N(clknet_leaf_19_clk),
    .D(net311),
    .RESET_B(net12),
    .SET_B(net266),
    .Q(net460));
 sky130_fd_sc_hd__dlrtn_1 c449 (.D(clknet_1_0__leaf_net452),
    .GATE_N(clknet_leaf_20_clk),
    .RESET_B(net828),
    .Q(net461));
 sky130_fd_sc_hd__dlymetal6s2s_1 c45 (.A(net21),
    .X(net23));
 sky130_fd_sc_hd__dfbbp_1 c450 (.CLK(clknet_leaf_18_clk),
    .D(net12),
    .RESET_B(clknet_1_0__leaf_net333),
    .SET_B(net811),
    .Q(net462));
 sky130_fd_sc_hd__and3_1 c451 (.A(net124),
    .B(net53),
    .C(net458),
    .X(net463));
 sky130_fd_sc_hd__sdfxbp_1 c452 (.CLK(clknet_leaf_20_clk),
    .D(net24),
    .SCD(clknet_1_0__leaf_net784),
    .SCE(net12),
    .Q(net464));
 sky130_fd_sc_hd__and2_0 c453 (.A(net270),
    .B(clknet_1_0__leaf_net337),
    .X(net465));
 sky130_fd_sc_hd__and2_1 c454 (.A(net754),
    .B(net776),
    .X(net466));
 sky130_fd_sc_hd__and2_0 c455 (.A(net461),
    .B(net265),
    .X(net467));
 sky130_fd_sc_hd__sdfxbp_1 c456 (.CLK(clknet_leaf_20_clk),
    .D(net189),
    .SCD(clknet_1_0__leaf_net465),
    .SCE(net447),
    .Q(net468));
 sky130_fd_sc_hd__sdfxtp_1 c457 (.CLK(clknet_leaf_20_clk),
    .D(clknet_1_1__leaf_net387),
    .SCD(net51),
    .SCE(clknet_1_1__leaf_net465),
    .Q(net469));
 sky130_fd_sc_hd__and3_1 c458 (.A(net469),
    .B(net881),
    .C(net461),
    .X(net470));
 sky130_fd_sc_hd__and2_0 c459 (.A(net459),
    .B(clknet_1_1__leaf_net130),
    .X(net471));
 sky130_fd_sc_hd__clkbuf_2 c46 (.A(net774),
    .X(net24));
 sky130_fd_sc_hd__dlrtn_1 c460 (.D(net463),
    .GATE_N(clknet_leaf_18_clk),
    .RESET_B(net457),
    .Q(net472));
 sky130_fd_sc_hd__and2_0 c461 (.A(net467),
    .B(net472),
    .X(net473));
 sky130_fd_sc_hd__and3_1 c462 (.A(net195),
    .B(net201),
    .C(net46),
    .X(net792));
 sky130_fd_sc_hd__and3_1 c463 (.A(net804),
    .B(net418),
    .C(net764),
    .X(net474));
 sky130_fd_sc_hd__and3_1 c464 (.A(net389),
    .B(net471),
    .C(net783),
    .X(net475));
 sky130_fd_sc_hd__dlrtp_1 c465 (.D(net217),
    .GATE(clknet_leaf_28_clk),
    .RESET_B(net394),
    .Q(net476));
 sky130_fd_sc_hd__and3_1 c466 (.A(net314),
    .B(net474),
    .C(net219),
    .X(net477));
 sky130_fd_sc_hd__sdfxtp_1 c467 (.CLK(clknet_leaf_21_clk),
    .D(net422),
    .SCD(net22),
    .SCE(net456),
    .Q(net478));
 sky130_fd_sc_hd__sdfxtp_1 c468 (.CLK(clknet_leaf_19_clk),
    .D(net4),
    .SCD(net249),
    .SCE(clknet_1_0__leaf_net337),
    .Q(net479));
 sky130_fd_sc_hd__and3_1 c469 (.A(net295),
    .B(net348),
    .C(net34),
    .X(net480));
 sky130_fd_sc_hd__and2_1 c47 (.A(net769),
    .B(net23),
    .X(net25));
 sky130_fd_sc_hd__and3_1 c470 (.A(net380),
    .B(net809),
    .C(net222),
    .X(net481));
 sky130_fd_sc_hd__and3_1 c471 (.A(net862),
    .B(net468),
    .C(net388),
    .X(net482));
 sky130_fd_sc_hd__dlrtp_1 c472 (.D(net22),
    .GATE(clknet_leaf_12_clk),
    .RESET_B(net40),
    .Q(net483));
 sky130_fd_sc_hd__dfbbn_1 c473 (.CLK_N(clknet_leaf_14_clk),
    .D(net265),
    .RESET_B(net475),
    .SET_B(net37),
    .Q(net484));
 sky130_fd_sc_hd__and3_1 c474 (.A(net478),
    .B(net483),
    .C(net4),
    .X(net485));
 sky130_fd_sc_hd__dfbbn_1 c475 (.CLK_N(clknet_leaf_17_clk),
    .D(net480),
    .RESET_B(clknet_1_0__leaf_net150),
    .SET_B(net470),
    .Q(net486));
 sky130_fd_sc_hd__dfbbp_1 c476 (.CLK(clknet_leaf_20_clk),
    .D(net810),
    .RESET_B(net484),
    .SET_B(net214),
    .Q(net487));
 sky130_fd_sc_hd__mux4_2 c477 (.A0(net358),
    .A1(net356),
    .A2(net401),
    .A3(net121),
    .S0(net755),
    .S1(net759),
    .X(net785));
 sky130_fd_sc_hd__dlrtp_1 c478 (.D(net388),
    .GATE(clknet_leaf_3_clk),
    .RESET_B(net360),
    .Q(net488));
 sky130_fd_sc_hd__sdfxbp_1 c479 (.CLK(clknet_leaf_13_clk),
    .D(net214),
    .SCD(net853),
    .SCE(net772),
    .Q(net489));
 sky130_fd_sc_hd__dfxtp_2 c48 (.CLK(clknet_leaf_6_clk),
    .D(net25),
    .Q(net26));
 sky130_fd_sc_hd__and2_1 c480 (.A(net325),
    .B(net215),
    .X(net490));
 sky130_fd_sc_hd__and3_1 c481 (.A(net21),
    .B(net489),
    .C(net756),
    .X(net491));
 sky130_fd_sc_hd__sdfxbp_1 c482 (.CLK(clknet_leaf_3_clk),
    .D(net203),
    .SCD(net482),
    .SCE(net418),
    .Q(net492));
 sky130_fd_sc_hd__sdfbbn_1 c487 (.CLK_N(clknet_leaf_16_clk),
    .D(clknet_1_1__leaf_net229),
    .RESET_B(net760),
    .SCD(net799),
    .SCE(net783),
    .SET_B(net785),
    .Q(net493));
 sky130_fd_sc_hd__sdfxtp_1 c488 (.CLK(clknet_leaf_16_clk),
    .D(net493),
    .SCD(net806),
    .SCE(net379),
    .Q(net494));
 sky130_fd_sc_hd__sdfrtp_1 c489 (.CLK(clknet_leaf_15_clk),
    .D(clknet_1_1__leaf_net150),
    .RESET_B(net466),
    .SCD(net877),
    .SCE(net125),
    .Q(net495));
 sky130_fd_sc_hd__clkbuf_2 c49 (.A(net766),
    .X(net27));
 sky130_fd_sc_hd__and3_1 c490 (.A(net243),
    .B(net365),
    .C(clknet_1_1__leaf_net789),
    .X(net496));
 sky130_fd_sc_hd__and3_1 c491 (.A(net219),
    .B(clknet_1_1__leaf_net337),
    .C(net240),
    .X(net497));
 sky130_fd_sc_hd__a2111o_1 c492 (.A1(net240),
    .A2(net363),
    .B1(net43),
    .C1(net339),
    .D1(net756),
    .X(net498));
 sky130_fd_sc_hd__sdfrtp_1 c493 (.CLK(clknet_leaf_16_clk),
    .D(net496),
    .RESET_B(clknet_1_1__leaf_net333),
    .SCD(net796),
    .SCE(net783),
    .Q(net499));
 sky130_fd_sc_hd__sdfxtp_1 c494 (.CLK(clknet_leaf_11_clk),
    .D(net772),
    .SCD(net375),
    .SCE(net498),
    .Q(net500));
 sky130_fd_sc_hd__a2111o_1 c495 (.A1(net760),
    .A2(net366),
    .B1(net804),
    .C1(net43),
    .D1(net99),
    .X(net794));
 sky130_fd_sc_hd__sdfxtp_1 c496 (.CLK(clknet_leaf_17_clk),
    .D(net145),
    .SCD(net770),
    .SCE(clknet_1_1__leaf_net150),
    .Q(net501));
 sky130_fd_sc_hd__and3_1 c497 (.A(net251),
    .B(net500),
    .C(net497),
    .X(net502));
 sky130_fd_sc_hd__or4bb_1 c498 (.A(net194),
    .B(net486),
    .C_N(clknet_1_0__leaf_net797),
    .D_N(net783),
    .X(net503));
 sky130_fd_sc_hd__sdfsbp_1 c499 (.CLK(clknet_leaf_16_clk),
    .D(net416),
    .SCD(net502),
    .SCE(net852),
    .SET_B(net759),
    .Q(net504));
 sky130_fd_sc_hd__buf_2 c50 (.A(net24),
    .X(net28));
 sky130_fd_sc_hd__dfbbn_1 c500 (.CLK_N(clknet_leaf_10_clk),
    .D(net40),
    .RESET_B(net226),
    .SET_B(net477),
    .Q(net505));
 sky130_fd_sc_hd__sdfbbp_1 c501 (.CLK(clknet_leaf_16_clk),
    .D(net503),
    .RESET_B(net371),
    .SCD(net505),
    .SCE(net805),
    .SET_B(net770),
    .Q(net793));
 sky130_fd_sc_hd__and3_1 c502 (.A(net494),
    .B(net504),
    .C(net501),
    .X(net506));
 sky130_fd_sc_hd__or4bb_1 c503 (.A(net499),
    .B(net37),
    .C_N(net506),
    .D_N(net782));
 sky130_fd_sc_hd__edfxbp_1 c504 (.CLK(clknet_leaf_32_clk),
    .D(net767),
    .DE(net246),
    .Q(net507));
 sky130_fd_sc_hd__dlclkp_4 c505 (.CLK(clknet_leaf_0_clk),
    .GATE(net246),
    .GCLK(net508));
 sky130_fd_sc_hd__and2_1 c506 (.A(net117),
    .B(net385),
    .X(net509));
 sky130_fd_sc_hd__clkbuf_1 c507 (.A(net399),
    .X(net510));
 sky130_fd_sc_hd__and2_0 c508 (.A(net115),
    .B(clknet_1_0__leaf_net508),
    .X(net511));
 sky130_fd_sc_hd__dfbbn_1 c509 (.CLK_N(clknet_leaf_27_clk),
    .D(net394),
    .RESET_B(clknet_1_1__leaf_net511),
    .SET_B(net384),
    .Q(net513),
    .Q_N(net512));
 sky130_fd_sc_hd__and2_2 c51 (.A(net27),
    .B(net19),
    .X(net29));
 sky130_fd_sc_hd__and2_4 c510 (.A(net758),
    .B(net765),
    .X(net514));
 sky130_fd_sc_hd__edfxtp_1 c511 (.CLK(clknet_leaf_33_clk),
    .D(net132),
    .DE(net902),
    .Q(net515));
 sky130_fd_sc_hd__and2_1 c512 (.A(net509),
    .B(net399),
    .X(net516));
 sky130_fd_sc_hd__sdlclkp_1 c513 (.CLK(clknet_leaf_31_clk),
    .GATE(net762),
    .SCE(net516),
    .GCLK(net517));
 sky130_fd_sc_hd__buf_1 c514 (.A(clknet_1_0__leaf_net396),
    .X(net518));
 sky130_fd_sc_hd__buf_1 c515 (.A(clknet_1_0__leaf_net517),
    .X(net519));
 sky130_fd_sc_hd__buf_1 c516 (.A(net515),
    .X(net520));
 sky130_fd_sc_hd__and2_1 c517 (.A(net520),
    .B(net510),
    .X(net521));
 sky130_fd_sc_hd__and2_1 c518 (.A(net521),
    .B(net118),
    .X(net522));
 sky130_fd_sc_hd__and2_0 c519 (.A(clknet_1_1__leaf_net517),
    .B(clknet_1_0__leaf_net519),
    .X(net523));
 sky130_fd_sc_hd__buf_1 c52 (.A(net854),
    .X(net30));
 sky130_fd_sc_hd__sdlclkp_2 c520 (.CLK(clknet_leaf_26_clk),
    .GATE(clknet_1_0__leaf_net519),
    .SCE(net522),
    .GCLK(net524));
 sky130_fd_sc_hd__and2_0 c521 (.A(clknet_1_1__leaf_net523),
    .B(clknet_1_0__leaf_net519),
    .X(net525));
 sky130_fd_sc_hd__dfbbp_1 c522 (.CLK(clknet_leaf_32_clk),
    .D(net845),
    .RESET_B(clknet_1_0__leaf_net525),
    .SET_B(net399),
    .Q(net788),
    .Q_N(net526));
 sky130_fd_sc_hd__and3_1 c523 (.A(net386),
    .B(net889),
    .C(net521),
    .X(net798));
 sky130_fd_sc_hd__sdlclkp_4 c524 (.CLK(clknet_leaf_27_clk),
    .GATE(clknet_1_1__leaf_net525),
    .SCE(clknet_1_0__leaf_net523),
    .GCLK(net527));
 sky130_fd_sc_hd__and2_0 c525 (.A(net381),
    .B(net257),
    .X(net528));
 sky130_fd_sc_hd__dfrbp_1 c526 (.CLK(clknet_leaf_28_clk),
    .D(net144),
    .RESET_B(net812),
    .Q(net529));
 sky130_fd_sc_hd__and3_1 c527 (.A(clknet_1_0__leaf_net142),
    .B(net778),
    .C(net510),
    .X(net530));
 sky130_fd_sc_hd__and2_0 c528 (.A(net250),
    .B(net803),
    .X(net531));
 sky130_fd_sc_hd__and2_0 c529 (.A(clknet_1_0__leaf_net156),
    .B(net776),
    .X(net532));
 sky130_fd_sc_hd__clkbuf_2 c53 (.A(net761),
    .X(net31));
 sky130_fd_sc_hd__and2_0 c530 (.A(net138),
    .B(net283),
    .X(net533));
 sky130_fd_sc_hd__dfrbp_1 c531 (.CLK(clknet_leaf_22_clk),
    .D(clknet_1_0__leaf_net405),
    .RESET_B(clknet_1_1__leaf_net156),
    .Q(net535),
    .Q_N(net534));
 sky130_fd_sc_hd__and2_1 c532 (.A(net531),
    .B(net783),
    .X(net536));
 sky130_fd_sc_hd__and2_1 c533 (.A(net385),
    .B(net769),
    .X(net537));
 sky130_fd_sc_hd__sdfbbn_1 c534 (.CLK_N(clknet_leaf_29_clk),
    .D(net254),
    .RESET_B(net536),
    .SCD(net767),
    .SCE(net271),
    .SET_B(net840),
    .Q(net538));
 sky130_fd_sc_hd__dfrtn_1 c535 (.CLK_N(clknet_leaf_28_clk),
    .D(net248),
    .RESET_B(clknet_1_0__leaf_net511),
    .Q(net539));
 sky130_fd_sc_hd__dfrtp_1 c536 (.CLK(clknet_leaf_25_clk),
    .D(net528),
    .RESET_B(net838),
    .Q(net540));
 sky130_fd_sc_hd__dfrtp_1 c537 (.CLK(clknet_leaf_26_clk),
    .D(net522),
    .RESET_B(net815),
    .Q(net541));
 sky130_fd_sc_hd__and2_0 c538 (.A(net761),
    .B(net428),
    .X(net542));
 sky130_fd_sc_hd__and2_0 c539 (.A(net7),
    .B(net880),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_2 c54 (.A(net756),
    .X(net32));
 sky130_fd_sc_hd__and2_2 c540 (.A(net510),
    .B(net268),
    .X(net544));
 sky130_fd_sc_hd__and2_1 c541 (.A(net529),
    .B(net400),
    .X(net545));
 sky130_fd_sc_hd__dfrtp_1 c542 (.CLK(clknet_leaf_26_clk),
    .D(net543),
    .RESET_B(net850),
    .Q(net546));
 sky130_fd_sc_hd__and3_1 c543 (.A(net545),
    .B(net386),
    .C(net138),
    .X(net547));
 sky130_fd_sc_hd__mux4_1 c544 (.A0(net541),
    .A1(net534),
    .A2(net522),
    .A3(net545),
    .S0(clknet_1_0__leaf_net519),
    .S1(net544),
    .X(net548));
 sky130_fd_sc_hd__and2_0 c545 (.A(net546),
    .B(net767),
    .X(net549));
 sky130_fd_sc_hd__and2_1 c546 (.A(net427),
    .B(net28),
    .X(net550));
 sky130_fd_sc_hd__sdfxbp_1 c547 (.CLK(clknet_leaf_2_clk),
    .D(clknet_1_0__leaf_net511),
    .SCD(net386),
    .SCE(net132),
    .Q(net551));
 sky130_fd_sc_hd__sdfxbp_1 c548 (.CLK(clknet_leaf_2_clk),
    .D(net532),
    .SCD(net445),
    .SCE(net318),
    .Q(net553),
    .Q_N(net552));
 sky130_fd_sc_hd__sdfxtp_1 c549 (.CLK(clknet_leaf_28_clk),
    .D(net544),
    .SCD(net815),
    .SCE(net168),
    .Q(net554));
 sky130_fd_sc_hd__dlymetal6s2s_1 c55 (.A(net26),
    .X(net33));
 sky130_fd_sc_hd__dfsbp_1 c550 (.CLK(clknet_leaf_2_clk),
    .D(net168),
    .SET_B(net798),
    .Q(net556),
    .Q_N(net555));
 sky130_fd_sc_hd__sdfxtp_1 c551 (.CLK(clknet_leaf_21_clk),
    .D(net299),
    .SCD(clknet_1_1__leaf_net429),
    .SCE(net8),
    .Q(net557));
 sky130_fd_sc_hd__and3_1 c552 (.A(net7),
    .B(net318),
    .C(net284),
    .X(net558));
 sky130_fd_sc_hd__and3_1 c553 (.A(net304),
    .B(net554),
    .C(net557),
    .X(net559));
 sky130_fd_sc_hd__and3_1 c554 (.A(net778),
    .B(net411),
    .C(clknet_1_0__leaf_net519),
    .X(net560));
 sky130_fd_sc_hd__and3_1 c555 (.A(net559),
    .B(net554),
    .C(net514),
    .X(net561));
 sky130_fd_sc_hd__sdfxtp_1 c556 (.CLK(clknet_leaf_1_clk),
    .D(net770),
    .SCD(net550),
    .SCE(net764),
    .Q(net562));
 sky130_fd_sc_hd__and2_0 c557 (.A(clknet_1_1__leaf_net508),
    .B(net18),
    .X(net563));
 sky130_fd_sc_hd__dfbbn_1 c558 (.CLK_N(clknet_leaf_0_clk),
    .D(clknet_1_0__leaf_net308),
    .RESET_B(net426),
    .SET_B(net514),
    .Q(net565),
    .Q_N(net564));
 sky130_fd_sc_hd__dfbbn_1 c559 (.CLK_N(clknet_leaf_3_clk),
    .D(net446),
    .RESET_B(net551),
    .SET_B(net552),
    .Q(net566));
 sky130_fd_sc_hd__dfrbp_2 c56 (.CLK(clknet_leaf_6_clk),
    .D(net33),
    .RESET_B(net30),
    .Q(net35),
    .Q_N(net34));
 sky130_fd_sc_hd__and3_1 c560 (.A(net284),
    .B(net763),
    .C(net127),
    .X(net567));
 sky130_fd_sc_hd__and3_1 c561 (.A(net18),
    .B(net768),
    .C(net555),
    .X(net568));
 sky130_fd_sc_hd__and3_1 c562 (.A(net568),
    .B(net566),
    .C(clknet_1_1__leaf_net519),
    .X(net569));
 sky130_fd_sc_hd__dfbbp_1 c563 (.CLK(clknet_leaf_21_clk),
    .D(net547),
    .RESET_B(net168),
    .SET_B(net542),
    .Q(net571),
    .Q_N(net570));
 sky130_fd_sc_hd__sdfxbp_1 c564 (.CLK(clknet_leaf_19_clk),
    .D(clknet_1_0__leaf_net298),
    .SCD(net755),
    .SCE(net568),
    .Q(net572));
 sky130_fd_sc_hd__and3_1 c565 (.A(net561),
    .B(net271),
    .C(net381),
    .X(net573));
 sky130_fd_sc_hd__sdfxbp_1 c566 (.CLK(clknet_leaf_22_clk),
    .D(net573),
    .SCD(net7),
    .SCE(clknet_1_1__leaf_net569),
    .Q(net574));
 sky130_fd_sc_hd__and3_1 c567 (.A(net115),
    .B(net258),
    .C(clknet_1_0__leaf_net423),
    .X(net575));
 sky130_fd_sc_hd__and3_1 c568 (.A(net542),
    .B(clknet_1_0__leaf_net129),
    .C(net756),
    .X(net576));
 sky130_fd_sc_hd__dfsbp_1 c569 (.CLK(clknet_leaf_23_clk),
    .D(net558),
    .SET_B(net811),
    .Q(net578),
    .Q_N(net577));
 sky130_fd_sc_hd__and2_1 c57 (.A(net827),
    .B(net9),
    .X(net36));
 sky130_fd_sc_hd__and3_1 c570 (.A(net425),
    .B(net419),
    .C(net318),
    .X(net579));
 sky130_fd_sc_hd__dfstp_1 c571 (.CLK(clknet_leaf_19_clk),
    .D(net861),
    .SET_B(clknet_1_1__leaf_net784),
    .Q(net580));
 sky130_fd_sc_hd__sdfxtp_1 c572 (.CLK(clknet_leaf_21_clk),
    .D(net409),
    .SCD(net262),
    .SCE(net323),
    .Q(net581));
 sky130_fd_sc_hd__and2_1 c573 (.A(net404),
    .B(net176),
    .X(net582));
 sky130_fd_sc_hd__and3_1 c574 (.A(net464),
    .B(clknet_1_1__leaf_net519),
    .C(net581),
    .X(net583));
 sky130_fd_sc_hd__dfstp_1 c575 (.CLK(clknet_leaf_28_clk),
    .D(net533),
    .SET_B(net414),
    .Q(net584));
 sky130_fd_sc_hd__and3_1 c576 (.A(net262),
    .B(net45),
    .C(net764),
    .X(net585));
 sky130_fd_sc_hd__sdfxtp_1 c577 (.CLK(clknet_leaf_29_clk),
    .D(net576),
    .SCD(net864),
    .SCE(net445),
    .Q(net586));
 sky130_fd_sc_hd__and2_1 c578 (.A(net581),
    .B(net739),
    .X(net587));
 sky130_fd_sc_hd__and3_1 c579 (.A(net587),
    .B(net199),
    .C(net759),
    .X(net588));
 sky130_fd_sc_hd__dfrtn_1 c58 (.CLK_N(clknet_leaf_7_clk),
    .D(net30),
    .RESET_B(net32),
    .Q(net37));
 sky130_fd_sc_hd__and2_0 c580 (.A(net773),
    .B(net324),
    .X(net589));
 sky130_fd_sc_hd__and2_0 c581 (.A(net255),
    .B(net780),
    .X(net590));
 sky130_fd_sc_hd__and3_1 c582 (.A(net588),
    .B(net428),
    .C(net760),
    .X(net591));
 sky130_fd_sc_hd__sdfxtp_1 c583 (.CLK(clknet_leaf_28_clk),
    .D(net538),
    .SCD(net837),
    .SCE(net591),
    .Q(net592));
 sky130_fd_sc_hd__dfbbn_1 c584 (.CLK_N(clknet_leaf_20_clk),
    .D(net589),
    .RESET_B(clknet_1_1__leaf_net298),
    .SET_B(net587),
    .Q(net593));
 sky130_fd_sc_hd__and2_1 c585 (.A(net473),
    .B(net582),
    .X(net594));
 sky130_fd_sc_hd__and3_1 c586 (.A(net592),
    .B(net586),
    .C(clknet_1_0__leaf_net300),
    .X(net595));
 sky130_fd_sc_hd__dfbbn_1 c587 (.CLK_N(clknet_leaf_20_clk),
    .D(net323),
    .RESET_B(net847),
    .SET_B(net594),
    .Q(net596));
 sky130_fd_sc_hd__sdfsbp_1 c588 (.CLK(clknet_leaf_23_clk),
    .D(net447),
    .SCD(net222),
    .SCE(net413),
    .SET_B(net819),
    .Q(net597));
 sky130_fd_sc_hd__sdfstp_1 c589 (.CLK(clknet_leaf_21_clk),
    .D(net585),
    .SCD(net583),
    .SCE(clknet_1_0__leaf_net129),
    .SET_B(net394),
    .Q(net598));
 sky130_fd_sc_hd__dfrtp_2 c59 (.CLK(clknet_leaf_6_clk),
    .D(net36),
    .RESET_B(net823),
    .Q(net38));
 sky130_fd_sc_hd__or4bb_1 c590 (.A(net537),
    .B(net13),
    .C_N(net768),
    .D_N(net346),
    .X(net599));
 sky130_fd_sc_hd__or4bb_1 c591 (.A(net127),
    .B(net768),
    .C_N(net321),
    .D_N(net803),
    .X(net600));
 sky130_fd_sc_hd__or4bb_1 c592 (.A(net182),
    .B(clknet_1_0__leaf_net569),
    .C_N(net766),
    .D_N(net34),
    .X(net601));
 sky130_fd_sc_hd__sdfbbn_1 c593 (.CLK_N(clknet_leaf_13_clk),
    .D(net492),
    .RESET_B(net389),
    .SCD(net143),
    .SCE(clknet_1_0__leaf_net595),
    .SET_B(net738),
    .Q(net602));
 sky130_fd_sc_hd__sdfstp_1 c594 (.CLK(clknet_leaf_18_clk),
    .D(net453),
    .SCD(net907),
    .SCE(net759),
    .SET_B(clknet_1_0__leaf_net800),
    .Q(net603));
 sky130_fd_sc_hd__dfbbp_1 c595 (.CLK(clknet_leaf_19_clk),
    .D(net143),
    .RESET_B(net833),
    .SET_B(net46),
    .Q(net604));
 sky130_fd_sc_hd__sdfbbp_1 c596 (.CLK(clknet_leaf_28_clk),
    .D(net761),
    .RESET_B(net481),
    .SCD(net602),
    .SCE(net534),
    .SET_B(clknet_1_1__leaf_net575),
    .Q(net605));
 sky130_fd_sc_hd__sdfbbn_1 c597 (.CLK_N(clknet_leaf_20_clk),
    .D(net444),
    .RESET_B(net381),
    .SCD(net603),
    .SCE(net157),
    .SET_B(net339),
    .Q(net606));
 sky130_fd_sc_hd__sdfstp_1 c598 (.CLK(clknet_leaf_23_clk),
    .D(net860),
    .SCD(net591),
    .SCE(net410),
    .SET_B(net826),
    .Q(net607));
 sky130_fd_sc_hd__sdfbbn_1 c599 (.CLK_N(clknet_leaf_22_clk),
    .D(net487),
    .RESET_B(net357),
    .SCD(net249),
    .SCE(net570),
    .SET_B(net600),
    .Q(net608));
 sky130_fd_sc_hd__dfrtp_2 c60 (.CLK(clknet_leaf_6_clk),
    .D(net32),
    .RESET_B(net36),
    .Q(net39));
 sky130_fd_sc_hd__sedfxbp_1 c600 (.CLK(clknet_leaf_23_clk),
    .D(net346),
    .DE(net607),
    .SCD(net599),
    .SCE(net512),
    .Q(net609));
 sky130_fd_sc_hd__sedfxbp_2 c601 (.CLK(clknet_leaf_23_clk),
    .D(net249),
    .DE(net557),
    .SCD(net604),
    .SCE(net892),
    .Q(net611),
    .Q_N(net610));
 sky130_fd_sc_hd__sdfbbp_1 c602 (.CLK(clknet_leaf_23_clk),
    .D(net166),
    .RESET_B(net601),
    .SCD(net892),
    .SCE(net537),
    .SET_B(net610),
    .Q(net612));
 sky130_fd_sc_hd__sdfbbn_1 c603 (.CLK_N(clknet_leaf_18_clk),
    .D(net157),
    .RESET_B(net462),
    .SCD(net127),
    .SCE(net315),
    .SET_B(net346),
    .Q(net613));
 sky130_fd_sc_hd__or4bb_1 c604 (.A(net897),
    .B(net580),
    .C_N(net613),
    .D_N(net611),
    .X(net614));
 sky130_fd_sc_hd__sdfbbn_1 c605 (.CLK_N(clknet_leaf_19_clk),
    .D(net614),
    .RESET_B(net594),
    .SCD(net841),
    .SCE(net147),
    .SET_B(net804),
    .Q(net615));
 sky130_fd_sc_hd__sedfxtp_1 c606 (.CLK(clknet_leaf_23_clk),
    .D(net456),
    .DE(net121),
    .SCD(net600),
    .SCE(net610),
    .Q(net616));
 sky130_fd_sc_hd__sedfxtp_1 c607 (.CLK(clknet_leaf_19_clk),
    .D(net888),
    .DE(clknet_1_1__leaf_net595),
    .SCD(net490),
    .SCE(net615),
    .Q(net617));
 sky130_fd_sc_hd__sdfbbp_1 c608 (.CLK(clknet_leaf_19_clk),
    .D(net470),
    .RESET_B(net835),
    .SCD(net417),
    .SCE(net871),
    .SET_B(net455),
    .Q(net618));
 sky130_fd_sc_hd__dfrtp_2 c61 (.CLK(clknet_leaf_8_clk),
    .D(net874),
    .RESET_B(net10),
    .Q(net40));
 sky130_fd_sc_hd__and3_1 c62 (.A(net31),
    .B(net14),
    .C(net765),
    .X(net41));
 sky130_fd_sc_hd__buf_1 c63 (.A(net2),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 c630 (.A(net397),
    .X(net619));
 sky130_fd_sc_hd__and2_0 c631 (.A(net776),
    .B(clknet_1_1__leaf_net527),
    .X(net620));
 sky130_fd_sc_hd__buf_1 c632 (.A(clknet_1_0__leaf_net129),
    .X(net621));
 sky130_fd_sc_hd__and3_1 c633 (.A(net757),
    .B(net384),
    .C(net389),
    .X(net622));
 sky130_fd_sc_hd__and2_0 c634 (.A(net118),
    .B(net761),
    .X(net623));
 sky130_fd_sc_hd__and2_0 c635 (.A(net119),
    .B(net397),
    .X(net624));
 sky130_fd_sc_hd__and2_0 c636 (.A(net762),
    .B(net901),
    .X(net625));
 sky130_fd_sc_hd__and2_1 c637 (.A(net764),
    .B(net775),
    .X(net626));
 sky130_fd_sc_hd__and2_0 c638 (.A(clknet_1_0__leaf_net527),
    .B(net389),
    .X(net627));
 sky130_fd_sc_hd__sdfxbp_1 c639 (.CLK(clknet_leaf_26_clk),
    .D(net623),
    .SCD(net773),
    .SCE(clknet_1_1__leaf_net524),
    .Q(net628));
 sky130_fd_sc_hd__dfsbp_2 c64 (.CLK(clknet_leaf_6_clk),
    .D(net25),
    .SET_B(net825),
    .Q(net780),
    .Q_N(net43));
 sky130_fd_sc_hd__and2_0 c640 (.A(net624),
    .B(clknet_1_1__leaf_net627),
    .X(net629));
 sky130_fd_sc_hd__and2_0 c641 (.A(net868),
    .B(net624),
    .X(net630));
 sky130_fd_sc_hd__and2_1 c642 (.A(net628),
    .B(net384),
    .X(net631));
 sky130_fd_sc_hd__and2_0 c643 (.A(net124),
    .B(net619),
    .X(net632));
 sky130_fd_sc_hd__sdfxbp_1 c644 (.CLK(clknet_leaf_27_clk),
    .D(net630),
    .SCD(net868),
    .SCE(net622),
    .Q(net633));
 sky130_fd_sc_hd__or4bb_2 c645 (.A(net633),
    .B(net761),
    .C_N(net626),
    .D_N(net774),
    .X(net634));
 sky130_fd_sc_hd__dfstp_1 c646 (.CLK(clknet_leaf_32_clk),
    .D(clknet_1_1__leaf_net629),
    .SET_B(clknet_1_0__leaf_net524),
    .Q(net635));
 sky130_fd_sc_hd__dlrbn_1 c647 (.D(net516),
    .GATE_N(clknet_leaf_31_clk),
    .RESET_B(net625),
    .Q(net637),
    .Q_N(net636));
 sky130_fd_sc_hd__dlrbn_1 c648 (.D(net632),
    .GATE_N(clknet_leaf_32_clk),
    .RESET_B(net763),
    .Q(net638));
 sky130_fd_sc_hd__dlrbp_1 c649 (.D(net622),
    .GATE(clknet_leaf_31_clk),
    .RESET_B(clknet_1_0__leaf_net518),
    .Q(net640),
    .Q_N(net639));
 sky130_fd_sc_hd__buf_1 c65 (.A(net32),
    .X(net44));
 sky130_fd_sc_hd__sedfxtp_1 c650 (.CLK(clknet_leaf_32_clk),
    .D(net638),
    .DE(clknet_1_0__leaf_net629),
    .SCD(net635),
    .SCE(net634),
    .Q(net641));
 sky130_fd_sc_hd__and2_1 c651 (.A(net384),
    .B(net513),
    .X(net642));
 sky130_fd_sc_hd__sdfxtp_1 c652 (.CLK(clknet_leaf_31_clk),
    .D(net867),
    .SCD(net141),
    .SCE(net642),
    .Q(net643));
 sky130_fd_sc_hd__sdfbbn_1 c653 (.CLK_N(clknet_leaf_32_clk),
    .D(net619),
    .RESET_B(net412),
    .SCD(clknet_1_0__leaf_net621),
    .SCE(net634),
    .SET_B(net641),
    .Q(net645),
    .Q_N(net644));
 sky130_fd_sc_hd__and2_0 c654 (.A(net530),
    .B(net261),
    .X(net646));
 sky130_fd_sc_hd__sdfxtp_2 c655 (.CLK(clknet_leaf_0_clk),
    .D(net756),
    .SCD(net120),
    .SCE(net132),
    .Q(net647));
 sky130_fd_sc_hd__and2_0 c656 (.A(net626),
    .B(net274),
    .X(net648));
 sky130_fd_sc_hd__and3_1 c657 (.A(clknet_1_0__leaf_net524),
    .B(net274),
    .C(clknet_1_0__leaf_net620),
    .X(net649));
 sky130_fd_sc_hd__and3_1 c658 (.A(net762),
    .B(net803),
    .C(net741),
    .X(net650));
 sky130_fd_sc_hd__sdfxtp_1 c659 (.CLK(clknet_leaf_31_clk),
    .D(net646),
    .SCD(clknet_1_0__leaf_net396),
    .SCE(net645),
    .Q(net651));
 sky130_fd_sc_hd__dfxtp_2 c66 (.CLK(clknet_leaf_6_clk),
    .D(net30),
    .Q(net45));
 sky130_fd_sc_hd__and2_0 c660 (.A(clknet_1_0__leaf_net627),
    .B(clknet_1_0__leaf_net620),
    .X(net652));
 sky130_fd_sc_hd__and3_1 c661 (.A(net411),
    .B(net762),
    .C(net740),
    .X(net653));
 sky130_fd_sc_hd__dfbbn_1 c662 (.CLK_N(clknet_leaf_31_clk),
    .D(net631),
    .RESET_B(net544),
    .SET_B(net647),
    .Q(net655),
    .Q_N(net654));
 sky130_fd_sc_hd__and2_0 c663 (.A(net649),
    .B(net776),
    .X(net656));
 sky130_fd_sc_hd__dfbbn_2 c664 (.CLK_N(clknet_leaf_31_clk),
    .D(net549),
    .RESET_B(net642),
    .SET_B(net631),
    .Q(net658),
    .Q_N(net657));
 sky130_fd_sc_hd__and2_0 c665 (.A(net645),
    .B(clknet_1_0__leaf_net518),
    .X(net659));
 sky130_fd_sc_hd__and3_1 c666 (.A(net650),
    .B(net761),
    .C(net644),
    .X(net660));
 sky130_fd_sc_hd__dfbbp_1 c667 (.CLK(clknet_leaf_33_clk),
    .D(net851),
    .RESET_B(clknet_1_0__leaf_net652),
    .SET_B(net514),
    .Q(net661));
 sky130_fd_sc_hd__and3_1 c668 (.A(net659),
    .B(net764),
    .C(net647),
    .X(net662));
 sky130_fd_sc_hd__sdfbbn_1 c669 (.CLK_N(clknet_leaf_31_clk),
    .D(net662),
    .RESET_B(clknet_1_1__leaf_net652),
    .SCD(net635),
    .SCE(net654),
    .SET_B(net509),
    .Q(net663));
 sky130_fd_sc_hd__and2_4 c67 (.A(net0),
    .B(net43),
    .X(net46));
 sky130_fd_sc_hd__a2111o_1 c670 (.A1(net625),
    .A2(net268),
    .B1(net658),
    .C1(clknet_1_1__leaf_net518),
    .D1(net152),
    .X(net664));
 sky130_fd_sc_hd__dlrbp_1 c671 (.D(net540),
    .GATE(clknet_leaf_25_clk),
    .RESET_B(net664),
    .Q(net665));
 sky130_fd_sc_hd__sdfxbp_1 c672 (.CLK(clknet_leaf_30_clk),
    .D(net117),
    .SCD(net439),
    .SCE(clknet_1_1__leaf_net656),
    .Q(net666));
 sky130_fd_sc_hd__and2_0 c673 (.A(net16),
    .B(net259),
    .X(net667));
 sky130_fd_sc_hd__sdfxbp_1 c674 (.CLK(clknet_leaf_33_clk),
    .D(net400),
    .SCD(net13),
    .SCE(net550),
    .Q(net668));
 sky130_fd_sc_hd__a2111o_1 c675 (.A1(net634),
    .A2(net775),
    .B1(net639),
    .C1(net445),
    .D1(net647),
    .X(net669));
 sky130_fd_sc_hd__sdfrbp_1 c676 (.CLK(clknet_leaf_0_clk),
    .D(net550),
    .RESET_B(net807),
    .SCD(net564),
    .SCE(net126),
    .Q(net670));
 sky130_fd_sc_hd__sdfxtp_1 c677 (.CLK(clknet_leaf_30_clk),
    .D(net31),
    .SCD(clknet_1_0__leaf_net656),
    .SCE(net544),
    .Q(net671));
 sky130_fd_sc_hd__dlrtn_1 c678 (.D(clknet_1_0__leaf_net429),
    .GATE_N(clknet_leaf_2_clk),
    .RESET_B(net16),
    .Q(net672));
 sky130_fd_sc_hd__mux4_1 c679 (.A0(net769),
    .A1(net315),
    .A2(net655),
    .A3(net647),
    .S0(net657),
    .S1(net859),
    .X(net673));
 sky130_fd_sc_hd__dfsbp_1 c68 (.CLK(clknet_leaf_7_clk),
    .D(net41),
    .SET_B(net10),
    .Q(net48),
    .Q_N(net47));
 sky130_fd_sc_hd__sdfxtp_1 c680 (.CLK(clknet_leaf_30_clk),
    .D(net848),
    .SCD(net669),
    .SCE(clknet_1_0__leaf_net301),
    .Q(net674));
 sky130_fd_sc_hd__and2_1 c681 (.A(net8),
    .B(net440),
    .X(net675));
 sky130_fd_sc_hd__sdfxtp_1 c682 (.CLK(clknet_leaf_30_clk),
    .D(net859),
    .SCD(net653),
    .SCE(clknet_1_0__leaf_net656),
    .Q(net676));
 sky130_fd_sc_hd__and3_1 c683 (.A(net635),
    .B(net514),
    .C(net765),
    .X(net677));
 sky130_fd_sc_hd__dfbbn_1 c684 (.CLK_N(clknet_leaf_33_clk),
    .D(net439),
    .RESET_B(net667),
    .SET_B(net514),
    .Q(net678));
 sky130_fd_sc_hd__and3_1 c685 (.A(net677),
    .B(net678),
    .C(net636),
    .X(net679));
 sky130_fd_sc_hd__and3_1 c686 (.A(net663),
    .B(net859),
    .C(net734),
    .X(net680));
 sky130_fd_sc_hd__and3_1 c687 (.A(net560),
    .B(net20),
    .C(net8),
    .X(net681));
 sky130_fd_sc_hd__dfbbn_1 c688 (.CLK_N(clknet_leaf_33_clk),
    .D(clknet_1_0__leaf_net652),
    .RESET_B(net778),
    .SET_B(net774),
    .Q(net683),
    .Q_N(net682));
 sky130_fd_sc_hd__dlrtn_1 c689 (.D(clknet_1_1__leaf_net621),
    .GATE_N(clknet_leaf_32_clk),
    .RESET_B(net679),
    .Q(net684));
 sky130_fd_sc_hd__and2_2 c69 (.A(net3),
    .B(net41),
    .X(net49));
 sky130_fd_sc_hd__dfbbp_1 c690 (.CLK(clknet_leaf_31_clk),
    .D(net842),
    .RESET_B(net681),
    .SET_B(net658),
    .Q(net685));
 sky130_fd_sc_hd__and3_1 c691 (.A(net432),
    .B(net643),
    .C(clknet_1_0__leaf_net301),
    .X(net686));
 sky130_fd_sc_hd__sdfxbp_1 c692 (.CLK(clknet_leaf_30_clk),
    .D(net673),
    .SCD(net686),
    .SCE(net400),
    .Q(net687));
 sky130_fd_sc_hd__or4bb_1 c693 (.A(net152),
    .B(net63),
    .C_N(net166),
    .D_N(net553),
    .X(net688));
 sky130_fd_sc_hd__and3_1 c694 (.A(net661),
    .B(net676),
    .C(net668),
    .X(net689));
 sky130_fd_sc_hd__sdfbbp_1 c695 (.CLK(clknet_leaf_30_clk),
    .D(net579),
    .RESET_B(net680),
    .SCD(net13),
    .SCE(net636),
    .SET_B(net684),
    .Q(net690));
 sky130_fd_sc_hd__mux4_1 c696 (.A0(net37),
    .A1(clknet_1_1__leaf_net518),
    .A2(clknet_1_1__leaf_net301),
    .A3(net45),
    .S0(net266),
    .S1(net733),
    .X(net691));
 sky130_fd_sc_hd__sdfrbp_1 c697 (.CLK(clknet_leaf_27_clk),
    .D(clknet_1_0__leaf_net153),
    .RESET_B(net830),
    .SCD(net685),
    .SCE(net514),
    .Q(net692));
 sky130_fd_sc_hd__sdfrtn_1 c698 (.CLK_N(clknet_leaf_33_clk),
    .D(net126),
    .RESET_B(net818),
    .SCD(net16),
    .SCE(net734),
    .Q(net693));
 sky130_fd_sc_hd__or4bb_1 c699 (.A(net445),
    .B(net261),
    .C_N(net658),
    .D_N(net775),
    .X(net694));
 sky130_fd_sc_hd__and2_1 c70 (.A(net767),
    .B(net44),
    .X(net50));
 sky130_fd_sc_hd__or4bb_1 c700 (.A(net885),
    .B(net556),
    .C_N(net62),
    .D_N(net274),
    .X(net695));
 sky130_fd_sc_hd__a2111o_1 c701 (.A1(net274),
    .A2(net660),
    .B1(net584),
    .C1(net680),
    .D1(net13),
    .X(net696));
 sky130_fd_sc_hd__sdfrtp_1 c702 (.CLK(clknet_leaf_31_clk),
    .D(net775),
    .RESET_B(net658),
    .SCD(net878),
    .SCE(net412),
    .Q(net697));
 sky130_fd_sc_hd__sdfrtp_1 c703 (.CLK(clknet_leaf_1_clk),
    .D(net590),
    .RESET_B(net813),
    .SCD(net196),
    .SCE(net16),
    .Q(net698));
 sky130_fd_sc_hd__sdfrtp_1 c704 (.CLK(clknet_leaf_30_clk),
    .D(net536),
    .RESET_B(net565),
    .SCD(net696),
    .SCE(net776),
    .Q(net699));
 sky130_fd_sc_hd__sdfbbn_1 c705 (.CLK_N(clknet_leaf_33_clk),
    .D(net412),
    .RESET_B(net675),
    .SCD(net869),
    .SCE(net763),
    .SET_B(net128),
    .Q(net700));
 sky130_fd_sc_hd__sdfsbp_1 c706 (.CLK(clknet_leaf_1_clk),
    .D(net13),
    .SCD(net647),
    .SCE(net126),
    .SET_B(net320),
    .Q(net702),
    .Q_N(net701));
 sky130_fd_sc_hd__sdfbbn_1 c707 (.CLK_N(clknet_leaf_2_clk),
    .D(net196),
    .RESET_B(net139),
    .SCD(net166),
    .SCE(net701),
    .SET_B(net675),
    .Q(net704),
    .Q_N(net703));
 sky130_fd_sc_hd__or4bb_1 c708 (.A(net258),
    .B(net700),
    .C_N(net690),
    .D_N(net321),
    .X(net705));
 sky130_fd_sc_hd__sdfbbp_1 c709 (.CLK(clknet_leaf_33_clk),
    .D(net693),
    .RESET_B(net694),
    .SCD(net858),
    .SCE(net704),
    .SET_B(net46),
    .Q(net707),
    .Q_N(net706));
 sky130_fd_sc_hd__dfstp_1 c71 (.CLK(clknet_leaf_7_clk),
    .D(net49),
    .SET_B(net32),
    .Q(net51));
 sky130_fd_sc_hd__a2111o_1 c710 (.A1(net707),
    .A2(net141),
    .B1(net695),
    .C1(net647),
    .D1(net703),
    .X(net708));
 sky130_fd_sc_hd__sdfbbn_1 c711 (.CLK_N(clknet_leaf_30_clk),
    .D(net125),
    .RESET_B(net143),
    .SCD(net674),
    .SCE(net707),
    .SET_B(net898),
    .Q(net709));
 sky130_fd_sc_hd__sdfbbn_1 c712 (.CLK_N(clknet_leaf_2_clk),
    .D(net691),
    .RESET_B(net886),
    .SCD(net689),
    .SCE(net705),
    .SET_B(net898),
    .Q(net710));
 sky130_fd_sc_hd__sdfsbp_1 c713 (.CLK(clknet_leaf_2_clk),
    .D(net132),
    .SCD(net704),
    .SCE(net899),
    .SET_B(net824),
    .Q(net711));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(net455),
    .A1(net28),
    .A2(net687),
    .A3(net596),
    .S0(net147),
    .S1(net905),
    .X(net712));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net756),
    .A1(net401),
    .A2(net491),
    .A3(net485),
    .S0(net906),
    .S1(net91),
    .X(net713));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net670),
    .A1(net567),
    .A2(net778),
    .A3(clknet_1_0__leaf_net575),
    .S0(net775),
    .S1(net16),
    .X(net714));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net688),
    .A1(net35),
    .A2(net74),
    .A3(net684),
    .S0(net611),
    .S1(net872),
    .X(net715));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(net612),
    .A1(net514),
    .A2(net472),
    .A3(net609),
    .S0(net709),
    .S1(net567),
    .X(net716));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net765),
    .A1(net181),
    .A2(net710),
    .A3(net803),
    .S0(net780),
    .S1(net745),
    .X(net717));
 sky130_fd_sc_hd__and2_1 c72 (.A(net804),
    .B(net755),
    .X(net52));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(clknet_1_1__leaf_net423),
    .A1(net1),
    .A2(net765),
    .A3(net267),
    .S0(net606),
    .S1(net744),
    .X(net718));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net539),
    .A1(net315),
    .A2(net476),
    .A3(net128),
    .S0(net692),
    .S1(net765),
    .X(net719));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net535),
    .A1(net755),
    .A2(net711),
    .A3(net321),
    .S0(net716),
    .S1(net637),
    .X(net720));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net128),
    .A1(net347),
    .A2(net257),
    .A3(net1),
    .S0(net755),
    .S1(net884),
    .X(net721));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net563),
    .A1(net757),
    .A2(net77),
    .A3(net717),
    .S0(net718),
    .S1(net143),
    .X(net722));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net120),
    .A1(net759),
    .A2(net578),
    .A3(net13),
    .S0(net746),
    .S1(net747),
    .X(net723));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net513),
    .A1(net764),
    .A2(net766),
    .A3(net438),
    .S0(net520),
    .S1(net763),
    .X(net724));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net509),
    .A1(net224),
    .A2(net665),
    .A3(net618),
    .S0(net166),
    .S1(net723),
    .X(net725));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(clknet_1_0__leaf_net300),
    .A1(net448),
    .A2(net655),
    .A3(net605),
    .S0(net749),
    .S1(net750),
    .X(net726));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(net267),
    .A1(net91),
    .A2(net571),
    .A3(net320),
    .S0(net45),
    .S1(net748),
    .X(net727));
 sky130_fd_sc_hd__dfstp_1 c73 (.CLK(clknet_leaf_6_clk),
    .D(net36),
    .SET_B(net25),
    .Q(net53));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(clknet_1_1__leaf_net620),
    .A1(net46),
    .A2(net648),
    .A3(clknet_1_1__leaf_net449),
    .S0(net608),
    .S1(net751),
    .X(net728));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net637),
    .A1(net450),
    .A2(net402),
    .A3(net757),
    .S0(net752),
    .S1(net753));
 sky130_fd_sc_hd__dfstp_1 c74 (.CLK(clknet_leaf_9_clk),
    .D(net50),
    .SET_B(net1),
    .Q(net54));
 sky130_fd_sc_hd__dlrbn_1 c75 (.D(net46),
    .GATE_N(clknet_leaf_17_clk),
    .RESET_B(net49),
    .Q(net56),
    .Q_N(net55));
 sky130_fd_sc_hd__and2_1 c76 (.A(net28),
    .B(net52),
    .X(net57));
 sky130_fd_sc_hd__and2_0 c77 (.A(net831),
    .B(net27),
    .X(net58));
 sky130_fd_sc_hd__dlrbn_1 c78 (.D(net42),
    .GATE_N(clknet_leaf_10_clk),
    .RESET_B(net881),
    .Q(net60),
    .Q_N(net59));
 sky130_fd_sc_hd__and2_1 c79 (.A(net48),
    .B(net19),
    .X(net61));
 sky130_fd_sc_hd__sdfrbp_1 c80 (.CLK(clknet_leaf_7_clk),
    .D(net50),
    .RESET_B(net52),
    .SCD(net57),
    .SCE(net59),
    .Q(net63),
    .Q_N(net62));
 sky130_fd_sc_hd__and2_1 c81 (.A(net63),
    .B(net58),
    .X(net64));
 sky130_fd_sc_hd__sdfbbn_1 c82 (.CLK_N(clknet_leaf_9_clk),
    .D(net856),
    .RESET_B(net64),
    .SCD(net32),
    .SCE(net49),
    .SET_B(net50),
    .Q(net66),
    .Q_N(net65));
 sky130_fd_sc_hd__and2_1 c83 (.A(net61),
    .B(net58),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 c84 (.A(net9),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 c85 (.A(net774),
    .X(net69));
 sky130_fd_sc_hd__and2_1 c86 (.A(net761),
    .B(net65),
    .X(net70));
 sky130_fd_sc_hd__and2_0 c87 (.A(net804),
    .B(net66),
    .X(net71));
 sky130_fd_sc_hd__dlrbp_1 c88 (.D(net67),
    .GATE(clknet_leaf_10_clk),
    .RESET_B(net42),
    .Q(net73),
    .Q_N(net72));
 sky130_fd_sc_hd__and2_1 c89 (.A(net21),
    .B(net29),
    .X(net74));
 sky130_fd_sc_hd__buf_1 c90 (.A(net768),
    .X(net75));
 sky130_fd_sc_hd__and3_1 c91 (.A(net58),
    .B(net34),
    .C(net756),
    .X(net76));
 sky130_fd_sc_hd__and2_1 c92 (.A(net51),
    .B(net757),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 c93 (.A(net75),
    .X(net78));
 sky130_fd_sc_hd__and2_1 c94 (.A(net47),
    .B(net14),
    .X(net79));
 sky130_fd_sc_hd__dlrbp_1 c95 (.D(net74),
    .GATE(clknet_leaf_12_clk),
    .RESET_B(net774),
    .Q(net81),
    .Q_N(net80));
 sky130_fd_sc_hd__and2_1 c96 (.A(net77),
    .B(net3),
    .X(net82));
 sky130_fd_sc_hd__and2_1 c97 (.A(net69),
    .B(net778),
    .X(net83));
 sky130_fd_sc_hd__dlrtn_1 c98 (.D(net68),
    .GATE_N(clknet_leaf_15_clk),
    .RESET_B(net27),
    .Q(net84));
 sky130_fd_sc_hd__dfbbn_1 c99 (.CLK_N(clknet_leaf_10_clk),
    .D(net83),
    .RESET_B(net72),
    .SET_B(net42),
    .Q(net86),
    .Q_N(net85));
 sky130_fd_sc_hd__sdfstp_1 merge732 (.CLK(clknet_leaf_28_clk),
    .D(clknet_1_1__leaf_net398),
    .SCD(net380),
    .SCE(clknet_1_1__leaf_net393),
    .SET_B(clknet_1_0__leaf_net287),
    .Q(net729));
 sky130_fd_sc_hd__dlxbn_1 s733 (.D(net89),
    .GATE_N(clknet_leaf_17_clk),
    .Q(net731),
    .Q_N(net730));
 sky130_fd_sc_hd__dlxbn_1 s734 (.D(net98),
    .GATE_N(clknet_leaf_8_clk),
    .Q(net732));
 sky130_fd_sc_hd__dlxbp_1 s735 (.D(net131),
    .GATE(clknet_leaf_29_clk),
    .Q(net734),
    .Q_N(net733));
 sky130_fd_sc_hd__dlxtn_2 s736 (.D(net309),
    .GATE_N(clknet_leaf_4_clk),
    .Q(net735));
 sky130_fd_sc_hd__dlxtn_1 s737 (.D(net322),
    .GATE_N(clknet_leaf_20_clk),
    .Q(net736));
 sky130_fd_sc_hd__dlxtn_1 s738 (.D(net326),
    .GATE_N(clknet_leaf_14_clk),
    .Q(net737));
 sky130_fd_sc_hd__dlxtp_1 s739 (.D(net341),
    .GATE(clknet_leaf_13_clk),
    .Q(net738));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s740 (.D(net430),
    .SLEEP_B(clknet_leaf_20_clk),
    .Q(net739));
 sky130_fd_sc_hd__dfxbp_1 s741 (.CLK(clknet_leaf_32_clk),
    .D(net548),
    .Q(net741),
    .Q_N(net740));
 sky130_fd_sc_hd__dfxbp_1 s742 (.CLK(clknet_leaf_24_clk),
    .D(net712),
    .Q(net742));
 sky130_fd_sc_hd__dfxtp_1 s743 (.CLK(clknet_leaf_3_clk),
    .D(net713),
    .Q(net743));
 sky130_fd_sc_hd__dfxtp_1 s744 (.CLK(clknet_leaf_29_clk),
    .D(net714),
    .Q(net744));
 sky130_fd_sc_hd__dfxtp_1 s745 (.CLK(clknet_leaf_3_clk),
    .D(net715),
    .Q(net745));
 sky130_fd_sc_hd__dlclkp_1 s746 (.CLK(clknet_leaf_24_clk),
    .GATE(net719),
    .GCLK(net746));
 sky130_fd_sc_hd__dlclkp_2 s747 (.CLK(clknet_leaf_25_clk),
    .GATE(net720),
    .GCLK(net747));
 sky130_fd_sc_hd__dlclkp_4 s748 (.CLK(clknet_leaf_22_clk),
    .GATE(net721),
    .GCLK(net748));
 sky130_fd_sc_hd__dlxbn_1 s749 (.D(net722),
    .GATE_N(clknet_leaf_28_clk),
    .Q(net749));
 sky130_fd_sc_hd__dlxbn_1 s750 (.D(net724),
    .GATE_N(clknet_leaf_28_clk),
    .Q(net750));
 sky130_fd_sc_hd__dlxbp_1 s751 (.D(net725),
    .GATE(clknet_leaf_25_clk),
    .Q(net751));
 sky130_fd_sc_hd__dlxtn_1 s752 (.D(net726),
    .GATE_N(clknet_leaf_25_clk),
    .Q(net752));
 sky130_fd_sc_hd__dlxtn_2 s753 (.D(net727),
    .GATE_N(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dlxtn_1 s754 (.D(net728),
    .GATE_N(clknet_leaf_25_clk),
    .Q(net753));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_4 input1 (.A(in0),
    .X(net754));
 sky130_fd_sc_hd__clkbuf_8 input2 (.A(in1),
    .X(net755));
 sky130_fd_sc_hd__buf_4 input3 (.A(in10),
    .X(net756));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(in11),
    .X(net757));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(in12),
    .X(net758));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(in13),
    .X(net759));
 sky130_fd_sc_hd__buf_4 input7 (.A(in14),
    .X(net760));
 sky130_fd_sc_hd__buf_4 input8 (.A(in15),
    .X(net761));
 sky130_fd_sc_hd__buf_2 input9 (.A(in16),
    .X(net762));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(in17),
    .X(net763));
 sky130_fd_sc_hd__buf_4 input11 (.A(in18),
    .X(net764));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(in19),
    .X(net765));
 sky130_fd_sc_hd__buf_2 input13 (.A(in2),
    .X(net766));
 sky130_fd_sc_hd__buf_4 input14 (.A(in20),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(in21),
    .X(net768));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(in22),
    .X(net769));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(in23),
    .X(net770));
 sky130_fd_sc_hd__buf_2 input18 (.A(in24),
    .X(net771));
 sky130_fd_sc_hd__buf_2 input19 (.A(in3),
    .X(net772));
 sky130_fd_sc_hd__buf_4 input20 (.A(in4),
    .X(net773));
 sky130_fd_sc_hd__buf_4 input21 (.A(in5),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(in6),
    .X(net775));
 sky130_fd_sc_hd__clkbuf_4 input23 (.A(in7),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(in8),
    .X(net777));
 sky130_fd_sc_hd__clkbuf_4 input25 (.A(in9),
    .X(net778));
 sky130_fd_sc_hd__buf_2 output26 (.A(net779),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output27 (.A(net780),
    .X(out10));
 sky130_fd_sc_hd__clkbuf_4 output28 (.A(net781),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_4 output29 (.A(net782),
    .X(out12));
 sky130_fd_sc_hd__clkbuf_4 output30 (.A(net783),
    .X(out13));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(clknet_1_1__leaf_net784),
    .X(out14));
 sky130_fd_sc_hd__buf_8 output32 (.A(net805),
    .X(out15));
 sky130_fd_sc_hd__clkbuf_4 output33 (.A(net786),
    .X(out16));
 sky130_fd_sc_hd__clkbuf_4 output34 (.A(net787),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output35 (.A(net788),
    .X(out18));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(clknet_1_1__leaf_net789),
    .X(out19));
 sky130_fd_sc_hd__clkbuf_4 output37 (.A(net790),
    .X(out2));
 sky130_fd_sc_hd__clkbuf_4 output38 (.A(net791),
    .X(out20));
 sky130_fd_sc_hd__clkbuf_4 output39 (.A(net792),
    .X(out21));
 sky130_fd_sc_hd__clkbuf_4 output40 (.A(net793),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_1 output41 (.A(net794),
    .X(out23));
 sky130_fd_sc_hd__clkbuf_4 output42 (.A(net795),
    .X(out24));
 sky130_fd_sc_hd__clkbuf_4 output43 (.A(net796),
    .X(out3));
 sky130_fd_sc_hd__clkbuf_1 output44 (.A(clknet_1_1__leaf_net797),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output45 (.A(net798),
    .X(out5));
 sky130_fd_sc_hd__clkbuf_4 output46 (.A(net799),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_1 output47 (.A(clknet_1_1__leaf_net800),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_4 output48 (.A(net801),
    .X(out8));
 sky130_fd_sc_hd__clkbuf_4 output49 (.A(net802),
    .X(out9));
 sky130_fd_sc_hd__buf_4 fanout50 (.A(net777),
    .X(net803));
 sky130_fd_sc_hd__buf_2 fanout51 (.A(net777),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net527 (.A(net527),
    .X(clknet_0_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net527 (.A(clknet_0_net527),
    .X(clknet_1_0__leaf_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net527 (.A(clknet_0_net527),
    .X(clknet_1_1__leaf_net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net627 (.A(net627),
    .X(clknet_0_net627));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net627 (.A(clknet_0_net627),
    .X(clknet_1_0__leaf_net627));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net627 (.A(clknet_0_net627),
    .X(clknet_1_1__leaf_net627));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net652 (.A(net652),
    .X(clknet_0_net652));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net652 (.A(clknet_0_net652),
    .X(clknet_1_0__leaf_net652));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net652 (.A(clknet_0_net652),
    .X(clknet_1_1__leaf_net652));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net629 (.A(net629),
    .X(clknet_0_net629));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net629 (.A(clknet_0_net629),
    .X(clknet_1_0__leaf_net629));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net629 (.A(clknet_0_net629),
    .X(clknet_1_1__leaf_net629));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net620 (.A(net620),
    .X(clknet_0_net620));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net620 (.A(clknet_0_net620),
    .X(clknet_1_0__leaf_net620));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net620 (.A(clknet_0_net620),
    .X(clknet_1_1__leaf_net620));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net656 (.A(net656),
    .X(clknet_0_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net656 (.A(clknet_0_net656),
    .X(clknet_1_0__leaf_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net656 (.A(clknet_0_net656),
    .X(clknet_1_1__leaf_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net524 (.A(net524),
    .X(clknet_0_net524));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net524 (.A(clknet_0_net524),
    .X(clknet_1_0__leaf_net524));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net524 (.A(clknet_0_net524),
    .X(clknet_1_1__leaf_net524));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net517 (.A(net517),
    .X(clknet_0_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net517 (.A(clknet_0_net517),
    .X(clknet_1_0__leaf_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net517 (.A(clknet_0_net517),
    .X(clknet_1_1__leaf_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net523 (.A(net523),
    .X(clknet_0_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net523 (.A(clknet_0_net523),
    .X(clknet_1_0__leaf_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net523 (.A(clknet_0_net523),
    .X(clknet_1_1__leaf_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net525 (.A(net525),
    .X(clknet_0_net525));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net525 (.A(clknet_0_net525),
    .X(clknet_1_0__leaf_net525));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net525 (.A(clknet_0_net525),
    .X(clknet_1_1__leaf_net525));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net519 (.A(net519),
    .X(clknet_0_net519));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net519 (.A(clknet_0_net519),
    .X(clknet_1_0__leaf_net519));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net519 (.A(clknet_0_net519),
    .X(clknet_1_1__leaf_net519));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net569 (.A(net569),
    .X(clknet_0_net569));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net569 (.A(clknet_0_net569),
    .X(clknet_1_0__leaf_net569));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net569 (.A(clknet_0_net569),
    .X(clknet_1_1__leaf_net569));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net508 (.A(net508),
    .X(clknet_0_net508));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net508 (.A(clknet_0_net508),
    .X(clknet_1_0__leaf_net508));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net508 (.A(clknet_0_net508),
    .X(clknet_1_1__leaf_net508));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net511 (.A(net511),
    .X(clknet_0_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net511 (.A(clknet_0_net511),
    .X(clknet_1_0__leaf_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net511 (.A(clknet_0_net511),
    .X(clknet_1_1__leaf_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net396 (.A(net396),
    .X(clknet_0_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_0__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_1__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net518 (.A(net518),
    .X(clknet_0_net518));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net518 (.A(clknet_0_net518),
    .X(clknet_1_0__leaf_net518));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net518 (.A(clknet_0_net518),
    .X(clknet_1_1__leaf_net518));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net398 (.A(net398),
    .X(clknet_0_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_0__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_1__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net337 (.A(net337),
    .X(clknet_0_net337));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net337 (.A(clknet_0_net337),
    .X(clknet_1_0__leaf_net337));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net337 (.A(clknet_0_net337),
    .X(clknet_1_1__leaf_net337));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net465 (.A(net465),
    .X(clknet_0_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net465 (.A(clknet_0_net465),
    .X(clknet_1_0__leaf_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net465 (.A(clknet_0_net465),
    .X(clknet_1_1__leaf_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net800 (.A(net800),
    .X(clknet_0_net800));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net800 (.A(clknet_0_net800),
    .X(clknet_1_0__leaf_net800));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net800 (.A(clknet_0_net800),
    .X(clknet_1_1__leaf_net800));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net452 (.A(net452),
    .X(clknet_0_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net452 (.A(clknet_0_net452),
    .X(clknet_1_0__leaf_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net452 (.A(clknet_0_net452),
    .X(clknet_1_1__leaf_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net333 (.A(net333),
    .X(clknet_0_net333));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net333 (.A(clknet_0_net333),
    .X(clknet_1_0__leaf_net333));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net333 (.A(clknet_0_net333),
    .X(clknet_1_1__leaf_net333));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net797 (.A(net797),
    .X(clknet_0_net797));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net797 (.A(clknet_0_net797),
    .X(clknet_1_0__leaf_net797));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net797 (.A(clknet_0_net797),
    .X(clknet_1_1__leaf_net797));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net229 (.A(net229),
    .X(clknet_0_net229));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net229 (.A(clknet_0_net229),
    .X(clknet_1_0__leaf_net229));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net229 (.A(clknet_0_net229),
    .X(clknet_1_1__leaf_net229));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net221 (.A(net221),
    .X(clknet_0_net221));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net221 (.A(clknet_0_net221),
    .X(clknet_1_0__leaf_net221));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net221 (.A(clknet_0_net221),
    .X(clknet_1_1__leaf_net221));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net142 (.A(net142),
    .X(clknet_0_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net142 (.A(clknet_0_net142),
    .X(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net142 (.A(clknet_0_net142),
    .X(clknet_1_1__leaf_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net423 (.A(net423),
    .X(clknet_0_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net423 (.A(clknet_0_net423),
    .X(clknet_1_0__leaf_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net423 (.A(clknet_0_net423),
    .X(clknet_1_1__leaf_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net575 (.A(net575),
    .X(clknet_0_net575));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net575 (.A(clknet_0_net575),
    .X(clknet_1_0__leaf_net575));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net575 (.A(clknet_0_net575),
    .X(clknet_1_1__leaf_net575));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net272 (.A(net272),
    .X(clknet_0_net272));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net272 (.A(clknet_0_net272),
    .X(clknet_1_0__leaf_net272));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net272 (.A(clknet_0_net272),
    .X(clknet_1_1__leaf_net272));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net150 (.A(net150),
    .X(clknet_0_net150));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net150 (.A(clknet_0_net150),
    .X(clknet_1_0__leaf_net150));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net150 (.A(clknet_0_net150),
    .X(clknet_1_1__leaf_net150));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net140 (.A(net140),
    .X(clknet_0_net140));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net140 (.A(clknet_0_net140),
    .X(clknet_1_0__leaf_net140));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net140 (.A(clknet_0_net140),
    .X(clknet_1_1__leaf_net140));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net149 (.A(net149),
    .X(clknet_0_net149));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net149 (.A(clknet_0_net149),
    .X(clknet_1_0__leaf_net149));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net149 (.A(clknet_0_net149),
    .X(clknet_1_1__leaf_net149));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net301 (.A(net301),
    .X(clknet_0_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net301 (.A(clknet_0_net301),
    .X(clknet_1_0__leaf_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net301 (.A(clknet_0_net301),
    .X(clknet_1_1__leaf_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net429 (.A(net429),
    .X(clknet_0_net429));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net429 (.A(clknet_0_net429),
    .X(clknet_1_0__leaf_net429));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net429 (.A(clknet_0_net429),
    .X(clknet_1_1__leaf_net429));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net308 (.A(net308),
    .X(clknet_0_net308));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net308 (.A(clknet_0_net308),
    .X(clknet_1_0__leaf_net308));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net308 (.A(clknet_0_net308),
    .X(clknet_1_1__leaf_net308));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net300 (.A(net300),
    .X(clknet_0_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net300 (.A(clknet_0_net300),
    .X(clknet_1_0__leaf_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net300 (.A(clknet_0_net300),
    .X(clknet_1_1__leaf_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net595 (.A(net595),
    .X(clknet_0_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_0__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_1__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net449 (.A(net449),
    .X(clknet_0_net449));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net449 (.A(clknet_0_net449),
    .X(clknet_1_0__leaf_net449));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net449 (.A(clknet_0_net449),
    .X(clknet_1_1__leaf_net449));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net153 (.A(net153),
    .X(clknet_0_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net153 (.A(clknet_0_net153),
    .X(clknet_1_0__leaf_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net153 (.A(clknet_0_net153),
    .X(clknet_1_1__leaf_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net151 (.A(net151),
    .X(clknet_0_net151));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net151 (.A(clknet_0_net151),
    .X(clknet_1_0__leaf_net151));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net151 (.A(clknet_0_net151),
    .X(clknet_1_1__leaf_net151));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net306 (.A(net306),
    .X(clknet_0_net306));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net306 (.A(clknet_0_net306),
    .X(clknet_1_0__leaf_net306));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net306 (.A(clknet_0_net306),
    .X(clknet_1_1__leaf_net306));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net298 (.A(net298),
    .X(clknet_0_net298));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net298 (.A(clknet_0_net298),
    .X(clknet_1_0__leaf_net298));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net298 (.A(clknet_0_net298),
    .X(clknet_1_1__leaf_net298));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net784 (.A(net784),
    .X(clknet_0_net784));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net784 (.A(clknet_0_net784),
    .X(clknet_1_0__leaf_net784));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net784 (.A(clknet_0_net784),
    .X(clknet_1_1__leaf_net784));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net135 (.A(net135),
    .X(clknet_0_net135));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net135 (.A(clknet_0_net135),
    .X(clknet_1_0__leaf_net135));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net135 (.A(clknet_0_net135),
    .X(clknet_1_1__leaf_net135));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net277 (.A(net277),
    .X(clknet_0_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net277 (.A(clknet_0_net277),
    .X(clknet_1_0__leaf_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net277 (.A(clknet_0_net277),
    .X(clknet_1_1__leaf_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net334 (.A(net334),
    .X(clknet_0_net334));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net334 (.A(clknet_0_net334),
    .X(clknet_1_0__leaf_net334));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net334 (.A(clknet_0_net334),
    .X(clknet_1_1__leaf_net334));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net336 (.A(net336),
    .X(clknet_0_net336));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net336 (.A(clknet_0_net336),
    .X(clknet_1_0__leaf_net336));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net336 (.A(clknet_0_net336),
    .X(clknet_1_1__leaf_net336));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net335 (.A(net335),
    .X(clknet_0_net335));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net335 (.A(clknet_0_net335),
    .X(clknet_1_0__leaf_net335));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net335 (.A(clknet_0_net335),
    .X(clknet_1_1__leaf_net335));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net287 (.A(net287),
    .X(clknet_0_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net287 (.A(clknet_0_net287),
    .X(clknet_1_0__leaf_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net287 (.A(clknet_0_net287),
    .X(clknet_1_1__leaf_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net405 (.A(net405),
    .X(clknet_0_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net405 (.A(clknet_0_net405),
    .X(clknet_1_0__leaf_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net405 (.A(clknet_0_net405),
    .X(clknet_1_1__leaf_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net290 (.A(net290),
    .X(clknet_0_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net290 (.A(clknet_0_net290),
    .X(clknet_1_0__leaf_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net290 (.A(clknet_0_net290),
    .X(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net129 (.A(net129),
    .X(clknet_0_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net129 (.A(clknet_0_net129),
    .X(clknet_1_0__leaf_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net129 (.A(clknet_0_net129),
    .X(clknet_1_1__leaf_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net621 (.A(net621),
    .X(clknet_0_net621));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net621 (.A(clknet_0_net621),
    .X(clknet_1_0__leaf_net621));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net621 (.A(clknet_0_net621),
    .X(clknet_1_1__leaf_net621));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net130 (.A(net130),
    .X(clknet_0_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net130 (.A(clknet_0_net130),
    .X(clknet_1_0__leaf_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net130 (.A(clknet_0_net130),
    .X(clknet_1_1__leaf_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net387 (.A(net387),
    .X(clknet_0_net387));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net387 (.A(clknet_0_net387),
    .X(clknet_1_0__leaf_net387));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net387 (.A(clknet_0_net387),
    .X(clknet_1_1__leaf_net387));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net393 (.A(net393),
    .X(clknet_0_net393));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net393 (.A(clknet_0_net393),
    .X(clknet_1_0__leaf_net393));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net393 (.A(clknet_0_net393),
    .X(clknet_1_1__leaf_net393));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net789 (.A(net789),
    .X(clknet_0_net789));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net789 (.A(clknet_0_net789),
    .X(clknet_1_0__leaf_net789));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net789 (.A(clknet_0_net789),
    .X(clknet_1_1__leaf_net789));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net162 (.A(net162),
    .X(clknet_0_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net162 (.A(clknet_0_net162),
    .X(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net162 (.A(clknet_0_net162),
    .X(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net156 (.A(net156),
    .X(clknet_0_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net156 (.A(clknet_0_net156),
    .X(clknet_1_0__leaf_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net156 (.A(clknet_0_net156),
    .X(clknet_1_1__leaf_net156));
 sky130_fd_sc_hd__buf_6 rebuffer1 (.A(net785),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net343),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net406),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net67),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net160),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net177),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net454),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net407),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net553),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net242),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net535),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net152),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net26),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net682),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net577),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net165),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net167),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net259),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net754),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net706),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net39),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net266),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net35),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net451),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net90),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net408),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net773),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net342),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net479),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net734),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net572),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net239),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net390),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net409),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net737),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net283),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net187),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net640),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net200),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net201),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net507),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net216),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net593),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net666),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net264),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net544),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net515),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net495),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net488),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net29),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net288),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net60),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net173),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net698),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net671),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net574),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net271),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net292),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net403),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net562),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net211),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net133),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net641),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net395),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net683),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net134),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net617),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net743),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net96),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net38),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net207),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net256),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net376),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net651),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net304),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net541),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net54),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net45),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net353),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net742),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net672),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net708),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net95),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net616),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net526),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net253),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net729),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net598),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net311),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(net55),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net40),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net291),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(net460),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net657),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(net702),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(net184),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(net397),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(net397),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(net15),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(net110),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(net697),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(net699),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(net597),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(net125),
    .X(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_B (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c25_X (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_SCE (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_SET_B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c27_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_X (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_X (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_D_N (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_D (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_X (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_SCE (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_D (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_RESET_B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_D (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c39_RESET_B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_X (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_SET_B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_SCD (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_SCE (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_DE (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A3 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_X (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_SET_B (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_D (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_SET_B (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_GATE (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_D (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_X (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c643_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_S1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_X (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold104_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_D (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_SCE (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_Q (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_SCE (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_D (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_SCE (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_D (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_D (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_X (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_SCD (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_C (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_D_N (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_X (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_SET_B (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_RESET_B (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_SCE (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_X (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net129_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_GCLK (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A3 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_D (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_D1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_SCD (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_SCD (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_X (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_D (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_SCE (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_SCE (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_D (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_RESET_B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_SCE (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_SCE (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_X (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_C (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_X (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_RESET_B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_RESET_B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c652_SCD (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_SET_B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_RESET_B (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_D (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_SCD (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_RESET_B (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_X (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_D (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_RESET_B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_D (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_RESET_B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_X (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_D (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_SCD (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_RESET_B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_X (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_SET_B (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_C (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_X (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S0 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_SCE (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_RESET_B (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_D (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_DE (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_X (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net150_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_X (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold12_A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_D1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_Q (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_B (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_Q (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net156_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_X (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_D (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_SCE (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_SCE (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_SCE (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_RESET_B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_SET_B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_RESET_B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_X (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_SCE (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_SCD (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_RESET_B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_X (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold5_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_Q (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S0 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_SCD (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_C_N (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_D (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_Q (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_RESET_B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_D (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_SCE (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_X (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_Q (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_D (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_X (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_SCE (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_SET_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_X (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_D (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_SCD (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_X (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c39_D (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c27_X (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_Q (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_D (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_RESET_B (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_RESET_B (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_X (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_D (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_SET_B (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_X (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_D (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_X (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_C (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_B (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_SCD (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_X (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_D (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_SCD (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c44_X (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_SCE (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_RESET_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_DE (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_X (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c47_B (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c45_X (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_D (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c50_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c46_X (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_D (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_RESET_B (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_GATE (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_DE (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_RESET_B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_D (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_SCE (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_RESET_B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_RESET_B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_X (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_D (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_SCD (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_SCD (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_X (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_SCD (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_SCD (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_D (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_X (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_D (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_Q (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold13_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c55_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c48_Q (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_B (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_S1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_D (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_SCE (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_RESET_B (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_SET_B (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_D (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_X (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_D (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_B (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_Q (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold22_A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_S0 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_SET_B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_Q_N (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_C (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A0 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A3 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_Q (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_C (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_Q (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_RESET_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c51_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c49_X (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold57_A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_SCE (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_RESET_B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_Q (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_D_N (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c657_B (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_B (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_D_N (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_S1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_B (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_Q (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c50_X (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_SCE (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_D (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_SET_B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_SET_B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_D (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_RESET_B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_X (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_C (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_GATE (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_SCD (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_Q (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net298_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_X (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c44_B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c28_X (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_D (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold75_A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_Q (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_D (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c53_X (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_C (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold89_A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_D (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_S0 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_B (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_Q (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_SCE (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_SCE (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_SET_B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_C (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_Q (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_Q (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_C (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_SCE (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_X (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_SET_B (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_RESET_B (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_RESET_B (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A0 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_X (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_D_N (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_C_N (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_B (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A3 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_Q (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_D (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_SCE (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_B (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_SCD (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_X (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_SCE (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_X (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_SET_B (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_C1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_Q_N (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_D_N (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c56_Q_N (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_C (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_SET_B (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_D (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_D_N (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_X (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_RESET_B (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_Q (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A0 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_SET_B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_X (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c58_Q (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_SET_B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_S0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold70_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_Q (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_RESET_B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_S1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_SCD (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_B (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_X (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_D (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_C (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_B (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_X (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c638_B (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_C (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_RESET_B (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_X (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold21_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c60_Q (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_SET_B (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_D (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_RESET_B (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_SET_B (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_X (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold98_A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold97_A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_B (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_Q (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_SET_B (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_B (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_C (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_Q (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_C (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_D (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_X (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold91_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c61_Q (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_D (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_RESET_B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_SCE (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_D (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_B (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_B (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_X (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A1 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A2 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_X (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold34_A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_D (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_X (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_D (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_SCE (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c653_RESET_B (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_X (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_SCE (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_SET_B (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_D (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_X (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_D (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_X (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_SCE (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_B (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_Q (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_Q_N (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_C1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_B1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_D (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_SCD (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_X (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_C1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_SCE (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_SCD (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_C (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_X (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_D (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_SCE (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_B (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_X (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net449_A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_X (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold78_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A3 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_Q (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A0 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_SET_B (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_X (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_D (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_SET_B (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_X (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_SET_B (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_C (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_RESET_B (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_X (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_SCE (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_RESET_B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_D (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_X (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_D (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_SCD (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_X (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A0 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_SET_B (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_X (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_Q (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_SCD (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_SCE (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_Q_N (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A1 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_SCE (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_SET_B (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_B (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_SET_B (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_SET_B (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_C (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_X (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_X (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_Q (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_B (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_SET_B (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold77_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_Q (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold46_A (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_SCE (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_RESET_B (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_D (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_X (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_Q (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_B (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_SCE (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_X (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_D (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_X (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S0 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_D_N (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_Q (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_Q_N (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_C_N (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A0 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S1 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_Q (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_C1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_SCD (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A3 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_D1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_C (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_SET_B (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_Q (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A2 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_Q (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A3 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_SET_B (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_Q (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_Q (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_SCD (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c32_X (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_C (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_Q (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_s749_D (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_X (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_s736_Q (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_B (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_s737_Q (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_C (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S1 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_C (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_SCE (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c33_X (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c28_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_X (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_D (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_RESET_B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_s733_D (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_X (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c57_B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c35_B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_X (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_X (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold19_A (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c31_A (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_SET_B (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_D (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_D (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A3 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_S0 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A1 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_B (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_SCD (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S0 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_D (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_B (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_C (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A0 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_D (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_C (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c54_A (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_D1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_C (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c33_A (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_D (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_B (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A1 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_B (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_A (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c44_A (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_B (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_A (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_D (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_B (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_SCE (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_C (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_SET_B (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_C (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A1 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_RESET_B (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_D1 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_B (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_B (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_B (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c645_B (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_B (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_D (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c53_A (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_B (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_B (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_B (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c658_A (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_GATE (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_C (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_SCE (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c648_RESET_B (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_B (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c30_B (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_D (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_B (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_C (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_SCE (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_C (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S0 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A2 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A0 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_C (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_C (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_B (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A0 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_C_N (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c49_A (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_B (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_D (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_C (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_B (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_A (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_B (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_SCD (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_D (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_D (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_B (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_C_N (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_B (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A2 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_B (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A0 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_B (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c47_A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_B (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_SCE (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_D (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_SET_B (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_SCD (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c32_A (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c25_A (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_SCD (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_B (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_B (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c30_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_B (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_D (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_SCE (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A2 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold27_A (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c639_SCD (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_SET_B (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_RESET_B (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_SET_B (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c645_D_N (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c46_A (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_B (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_B (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S0 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_D (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_D_N (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A2 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_B (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A2 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_SCE (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_B (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_B (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_B (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_RESET_B (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_B (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_B1 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_output27_A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_Q (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_B (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_output29_A (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_D_N (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_Q (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_output30_A (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_B (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_D_N (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_SCE (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_SCE (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_C (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_SCE (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_X (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net784_A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_X (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_output37_A (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_SCD (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_SCE (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_X (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_output43_A (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_SCD (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_SCD (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_X (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_SET_B (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_X (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_output49_A (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_B (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_SCD (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_RESET_B (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_RESET_B (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_X (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_X (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_A (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_SCE (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_C (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A3 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c658_B (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_D_N (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_S1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_X (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_SET_B (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_B1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_CLK_N (.DIODE(clknet_leaf_28_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_CLK (.DIODE(clknet_leaf_28_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_CLK (.DIODE(clknet_leaf_28_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_CLK (.DIODE(clknet_leaf_28_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge732_CLK (.DIODE(clknet_leaf_28_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_CLK (.DIODE(clknet_leaf_28_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s749_GATE_N (.DIODE(clknet_leaf_28_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s750_GATE_N (.DIODE(clknet_leaf_28_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_CLK (.DIODE(clknet_leaf_28_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_GATE (.DIODE(clknet_leaf_28_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_X (.DIODE(clknet_leaf_28_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_X (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_X (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_X (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_X (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_B (.DIODE(clknet_1_0__leaf_net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_GATE (.DIODE(clknet_1_0__leaf_net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_B (.DIODE(clknet_1_0__leaf_net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S0 (.DIODE(clknet_1_0__leaf_net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_C (.DIODE(clknet_1_0__leaf_net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net519_X (.DIODE(clknet_1_0__leaf_net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_D (.DIODE(clknet_1_0__leaf_net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_B (.DIODE(clknet_1_0__leaf_net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_C (.DIODE(clknet_1_0__leaf_net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_SET_B (.DIODE(clknet_1_0__leaf_net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net800_X (.DIODE(clknet_1_0__leaf_net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_RESET_B (.DIODE(clknet_1_0__leaf_net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_RESET_B (.DIODE(clknet_1_0__leaf_net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net150_X (.DIODE(clknet_1_0__leaf_net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_B (.DIODE(clknet_1_0__leaf_net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_C (.DIODE(clknet_1_0__leaf_net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A0 (.DIODE(clknet_1_0__leaf_net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net300_X (.DIODE(clknet_1_0__leaf_net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_SCE (.DIODE(clknet_1_1__leaf_net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_SCE (.DIODE(clknet_1_1__leaf_net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_SCE (.DIODE(clknet_1_1__leaf_net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net300_X (.DIODE(clknet_1_1__leaf_net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net153_A (.DIODE(clknet_0_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net153_A (.DIODE(clknet_0_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net153_X (.DIODE(clknet_0_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_RESET_B (.DIODE(clknet_1_0__leaf_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_D (.DIODE(clknet_1_0__leaf_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net153_X (.DIODE(clknet_1_0__leaf_net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_RESET_B (.DIODE(clknet_1_0__leaf_net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_SCD (.DIODE(clknet_1_0__leaf_net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net784_X (.DIODE(clknet_1_0__leaf_net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_SET_B (.DIODE(clknet_1_1__leaf_net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_output31_A (.DIODE(clknet_1_1__leaf_net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net784_X (.DIODE(clknet_1_1__leaf_net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A (.DIODE(clknet_1_0__leaf_net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_B (.DIODE(clknet_1_0__leaf_net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net135_X (.DIODE(clknet_1_0__leaf_net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net129_A (.DIODE(clknet_0_net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net129_A (.DIODE(clknet_0_net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net129_X (.DIODE(clknet_0_net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_B (.DIODE(clknet_1_0__leaf_net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_SCE (.DIODE(clknet_1_0__leaf_net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A (.DIODE(clknet_1_0__leaf_net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net129_X (.DIODE(clknet_1_0__leaf_net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B (.DIODE(clknet_1_1__leaf_net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A (.DIODE(clknet_1_1__leaf_net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_SCE (.DIODE(clknet_1_1__leaf_net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net129_X (.DIODE(clknet_1_1__leaf_net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_SCD (.DIODE(clknet_1_0__leaf_net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B (.DIODE(clknet_1_0__leaf_net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_B (.DIODE(clknet_1_0__leaf_net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net130_X (.DIODE(clknet_1_0__leaf_net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_B (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_D (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_B (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold5_X (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_RESET_B (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_RESET_B (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold13_X (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_SET_B (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_D (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold21_X (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_A (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_RESET_B (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold27_X (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_SCD (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_D (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_C (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold33_X (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold72_X (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_RESET_B (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_B (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold77_X (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net582));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
