module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net644;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net752;
 wire clknet_1_0__leaf_net752;
 wire clknet_1_1__leaf_net752;
 wire clknet_0_net751;
 wire clknet_1_0__leaf_net751;
 wire clknet_1_1__leaf_net751;
 wire clknet_0_net596;
 wire clknet_1_0__leaf_net596;
 wire clknet_1_1__leaf_net596;
 wire clknet_0_net750;
 wire clknet_1_0__leaf_net750;
 wire clknet_1_1__leaf_net750;
 wire clknet_0_net617;
 wire clknet_1_0__leaf_net617;
 wire clknet_1_1__leaf_net617;
 wire clknet_0_net695;
 wire clknet_1_0__leaf_net695;
 wire clknet_1_1__leaf_net695;
 wire clknet_0_net735;
 wire clknet_1_0__leaf_net735;
 wire clknet_1_1__leaf_net735;
 wire clknet_0_net734;
 wire clknet_1_0__leaf_net734;
 wire clknet_1_1__leaf_net734;
 wire clknet_0_net694;
 wire clknet_1_0__leaf_net694;
 wire clknet_1_1__leaf_net694;
 wire clknet_0_net582;
 wire clknet_1_0__leaf_net582;
 wire clknet_1_1__leaf_net582;
 wire clknet_0_net471;
 wire clknet_1_0__leaf_net471;
 wire clknet_1_1__leaf_net471;
 wire clknet_0_net472;
 wire clknet_1_0__leaf_net472;
 wire clknet_1_1__leaf_net472;
 wire clknet_0_net733;
 wire clknet_1_0__leaf_net733;
 wire clknet_1_1__leaf_net733;
 wire clknet_0_net448;
 wire clknet_1_0__leaf_net448;
 wire clknet_1_1__leaf_net448;
 wire clknet_0_net485;
 wire clknet_1_0__leaf_net485;
 wire clknet_1_1__leaf_net485;
 wire clknet_0_net438;
 wire clknet_1_0__leaf_net438;
 wire clknet_1_1__leaf_net438;
 wire clknet_0_net577;
 wire clknet_1_0__leaf_net577;
 wire clknet_1_1__leaf_net577;
 wire clknet_0_net548;
 wire clknet_1_0__leaf_net548;
 wire clknet_1_1__leaf_net548;
 wire clknet_0_net437;
 wire clknet_1_0__leaf_net437;
 wire clknet_1_1__leaf_net437;
 wire clknet_0_net455;
 wire clknet_1_0__leaf_net455;
 wire clknet_1_1__leaf_net455;
 wire clknet_0_net478;
 wire clknet_1_0__leaf_net478;
 wire clknet_1_1__leaf_net478;
 wire clknet_0_net443;
 wire clknet_1_0__leaf_net443;
 wire clknet_1_1__leaf_net443;
 wire clknet_0_net439;
 wire clknet_1_0__leaf_net439;
 wire clknet_1_1__leaf_net439;
 wire clknet_0_net545;
 wire clknet_1_0__leaf_net545;
 wire clknet_1_1__leaf_net545;
 wire clknet_0_net440;
 wire clknet_1_0__leaf_net440;
 wire clknet_1_1__leaf_net440;
 wire clknet_0_net863;
 wire clknet_1_0__leaf_net863;
 wire clknet_1_1__leaf_net863;
 wire clknet_0_net292;
 wire clknet_1_0__leaf_net292;
 wire clknet_1_1__leaf_net292;
 wire clknet_0_net290;
 wire clknet_1_0__leaf_net290;
 wire clknet_1_1__leaf_net290;
 wire clknet_0_net716;
 wire clknet_1_0__leaf_net716;
 wire clknet_1_1__leaf_net716;
 wire clknet_0_net249;
 wire clknet_1_0__leaf_net249;
 wire clknet_1_1__leaf_net249;
 wire clknet_0_net266;
 wire clknet_1_0__leaf_net266;
 wire clknet_1_1__leaf_net266;
 wire clknet_0_net270;
 wire clknet_1_0__leaf_net270;
 wire clknet_1_1__leaf_net270;
 wire clknet_0_net387;
 wire clknet_1_0__leaf_net387;
 wire clknet_1_1__leaf_net387;
 wire clknet_0_net269;
 wire clknet_1_0__leaf_net269;
 wire clknet_1_1__leaf_net269;
 wire clknet_0_net715;
 wire clknet_1_0__leaf_net715;
 wire clknet_1_1__leaf_net715;
 wire clknet_0_net251;
 wire clknet_1_0__leaf_net251;
 wire clknet_1_1__leaf_net251;
 wire clknet_0_net693;
 wire clknet_1_0__leaf_net693;
 wire clknet_1_1__leaf_net693;
 wire clknet_0_net237;
 wire clknet_1_0__leaf_net237;
 wire clknet_1_1__leaf_net237;
 wire clknet_0_net241;
 wire clknet_1_0__leaf_net241;
 wire clknet_1_1__leaf_net241;
 wire clknet_0_net121;
 wire clknet_1_0__leaf_net121;
 wire clknet_1_1__leaf_net121;
 wire clknet_0_net230;
 wire clknet_1_0__leaf_net230;
 wire clknet_1_1__leaf_net230;
 wire clknet_0_net357;
 wire clknet_1_0__leaf_net357;
 wire clknet_1_1__leaf_net357;
 wire clknet_0_net360;
 wire clknet_1_0__leaf_net360;
 wire clknet_1_1__leaf_net360;
 wire clknet_0_net366;
 wire clknet_1_0__leaf_net366;
 wire clknet_1_1__leaf_net366;
 wire clknet_0_net232;
 wire clknet_1_0__leaf_net232;
 wire clknet_1_1__leaf_net232;
 wire clknet_0_net890;
 wire clknet_1_0__leaf_net890;
 wire clknet_1_1__leaf_net890;
 wire clknet_0_net233;
 wire clknet_1_0__leaf_net233;
 wire clknet_1_1__leaf_net233;
 wire clknet_0_net117;
 wire clknet_1_0__leaf_net117;
 wire clknet_1_1__leaf_net117;
 wire clknet_0_net469;
 wire clknet_1_0__leaf_net469;
 wire clknet_1_1__leaf_net469;
 wire clknet_0_net124;
 wire clknet_1_0__leaf_net124;
 wire clknet_1_1__leaf_net124;
 wire clknet_0_net118;
 wire clknet_1_0__leaf_net118;
 wire clknet_1_1__leaf_net118;
 wire clknet_0_net132;
 wire clknet_1_0__leaf_net132;
 wire clknet_1_1__leaf_net132;
 wire clknet_0_net140;
 wire clknet_1_0__leaf_net140;
 wire clknet_1_1__leaf_net140;
 wire clknet_0_net866;
 wire clknet_1_0__leaf_net866;
 wire clknet_1_1__leaf_net866;
 wire clknet_0_net412;
 wire clknet_1_0__leaf_net412;
 wire clknet_1_1__leaf_net412;
 wire clknet_0_net144;
 wire clknet_1_0__leaf_net144;
 wire clknet_1_1__leaf_net144;
 wire clknet_0_net143;
 wire clknet_1_0__leaf_net143;
 wire clknet_1_1__leaf_net143;
 wire clknet_0_net142;
 wire clknet_1_0__leaf_net142;
 wire clknet_1_1__leaf_net142;
 wire clknet_0_net493;
 wire clknet_1_0__leaf_net493;
 wire clknet_1_1__leaf_net493;
 wire clknet_0_net282;
 wire clknet_1_0__leaf_net282;
 wire clknet_1_1__leaf_net282;
 wire clknet_0_net149;
 wire clknet_1_0__leaf_net149;
 wire clknet_1_1__leaf_net149;
 wire clknet_0_net134;
 wire clknet_1_0__leaf_net134;
 wire clknet_1_1__leaf_net134;
 wire clknet_0_net137;
 wire clknet_1_0__leaf_net137;
 wire clknet_1_1__leaf_net137;
 wire clknet_0_net263;
 wire clknet_1_0__leaf_net263;
 wire clknet_1_1__leaf_net263;
 wire clknet_0_net268;
 wire clknet_1_0__leaf_net268;
 wire clknet_1_1__leaf_net268;
 wire clknet_0_net489;
 wire clknet_1_0__leaf_net489;
 wire clknet_1_1__leaf_net489;
 wire clknet_0_net383;
 wire clknet_1_0__leaf_net383;
 wire clknet_1_1__leaf_net383;
 wire clknet_0_net386;
 wire clknet_1_0__leaf_net386;
 wire clknet_1_1__leaf_net386;
 wire clknet_0_net382;
 wire clknet_1_0__leaf_net382;
 wire clknet_1_1__leaf_net382;
 wire clknet_0_net376;
 wire clknet_1_0__leaf_net376;
 wire clknet_1_1__leaf_net376;
 wire clknet_0_net129;
 wire clknet_1_0__leaf_net129;
 wire clknet_1_1__leaf_net129;
 wire clknet_0_net139;
 wire clknet_1_0__leaf_net139;
 wire clknet_1_1__leaf_net139;
 wire clknet_0_net120;
 wire clknet_1_0__leaf_net120;
 wire clknet_1_1__leaf_net120;
 wire clknet_0_net463;
 wire clknet_1_0__leaf_net463;
 wire clknet_1_1__leaf_net463;
 wire clknet_0_net515;
 wire clknet_1_0__leaf_net515;
 wire clknet_1_1__leaf_net515;
 wire clknet_0_net122;
 wire clknet_1_0__leaf_net122;
 wire clknet_1_1__leaf_net122;
 wire clknet_0_net597;
 wire clknet_1_0__leaf_net597;
 wire clknet_1_1__leaf_net597;
 wire clknet_0_net127;
 wire clknet_1_0__leaf_net127;
 wire clknet_1_1__leaf_net127;
 wire clknet_0_net125;
 wire clknet_1_0__leaf_net125;
 wire clknet_1_1__leaf_net125;
 wire clknet_0_net116;
 wire clknet_1_0__leaf_net116;
 wire clknet_1_1__leaf_net116;
 wire clknet_0_net468;
 wire clknet_1_0__leaf_net468;
 wire clknet_1_1__leaf_net468;
 wire clknet_0_net465;
 wire clknet_1_0__leaf_net465;
 wire clknet_1_1__leaf_net465;
 wire clknet_0_net619;
 wire clknet_1_0__leaf_net619;
 wire clknet_1_1__leaf_net619;
 wire clknet_0_net572;
 wire clknet_1_0__leaf_net572;
 wire clknet_1_1__leaf_net572;
 wire clknet_0_net112;
 wire clknet_1_0__leaf_net112;
 wire clknet_1_1__leaf_net112;
 wire clknet_0_net114;
 wire clknet_1_0__leaf_net114;
 wire clknet_1_1__leaf_net114;
 wire clknet_0_net107;
 wire clknet_1_0__leaf_net107;
 wire clknet_1_1__leaf_net107;
 wire clknet_0_net113;
 wire clknet_1_0__leaf_net113;
 wire clknet_1_1__leaf_net113;
 wire clknet_0_net239;
 wire clknet_1_0__leaf_net239;
 wire clknet_1_1__leaf_net239;
 wire clknet_0_net592;
 wire clknet_1_0__leaf_net592;
 wire clknet_1_1__leaf_net592;
 wire clknet_0_net457;
 wire clknet_1_0__leaf_net457;
 wire clknet_1_1__leaf_net457;
 wire clknet_0_net119;
 wire clknet_1_0__leaf_net119;
 wire clknet_1_1__leaf_net119;
 wire clknet_0_net126;
 wire clknet_1_0__leaf_net126;
 wire clknet_1_1__leaf_net126;
 wire clknet_0_net884;
 wire clknet_1_0__leaf_net884;
 wire clknet_1_1__leaf_net884;
 wire clknet_0_net170;
 wire clknet_1_0__leaf_net170;
 wire clknet_1_1__leaf_net170;
 wire clknet_0_net136;
 wire clknet_1_0__leaf_net136;
 wire clknet_1_1__leaf_net136;
 wire clknet_0_net103;
 wire clknet_1_0__leaf_net103;
 wire clknet_1_1__leaf_net103;
 wire clknet_0_net550;
 wire clknet_1_0__leaf_net550;
 wire clknet_1_1__leaf_net550;
 wire clknet_0_net560;
 wire clknet_1_0__leaf_net560;
 wire clknet_1_1__leaf_net560;
 wire clknet_0_net551;
 wire clknet_1_0__leaf_net551;
 wire clknet_1_1__leaf_net551;
 wire clknet_0_net350;
 wire clknet_1_0__leaf_net350;
 wire clknet_1_1__leaf_net350;
 wire clknet_0_net354;
 wire clknet_1_0__leaf_net354;
 wire clknet_1_1__leaf_net354;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net989;
 wire net990;
 wire net991;
 wire net993;
 wire net995;
 wire net960;
 wire net988;
 wire net992;
 wire net994;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;

 sky130_fd_sc_hd__xnor2_2 c100 (.A(net24),
    .B(net22),
    .Y(net32));
 sky130_fd_sc_hd__a41o_2 c101 (.A1(net7),
    .A2(net4),
    .A3(net31),
    .A4(net26),
    .B1(net29),
    .X(net33));
 sky130_fd_sc_hd__xnor2_2 c102 (.A(net33),
    .B(net860),
    .Y(net34));
 sky130_fd_sc_hd__a21bo_1 c103 (.A1(net26),
    .A2(net29),
    .B1_N(net860),
    .X(net35));
 sky130_fd_sc_hd__sdfrbp_1 c104 (.CLK(clknet_4_4_0_clk),
    .D(net807),
    .RESET_B(net987),
    .SCD(net34),
    .SCE(net922),
    .Q(net37),
    .Q_N(net36));
 sky130_fd_sc_hd__xnor2_4 c105 (.A(net23),
    .B(net27),
    .Y(net38));
 sky130_fd_sc_hd__a21bo_1 c106 (.A1(net37),
    .A2(net35),
    .B1_N(net915),
    .X(net39));
 sky130_fd_sc_hd__a21bo_1 c107 (.A1(net31),
    .A2(net30),
    .B1_N(net39),
    .X(net40));
 sky130_fd_sc_hd__a21bo_2 c108 (.A1(net39),
    .A2(net800),
    .B1_N(net837),
    .X(net41));
 sky130_fd_sc_hd__mux4_1 c109 (.A0(net40),
    .A1(net24),
    .A2(net904),
    .A3(net22),
    .S0(net41),
    .S1(net38),
    .X(net42));
 sky130_fd_sc_hd__sdfrbp_2 c110 (.CLK(clknet_4_4_0_clk),
    .D(net806),
    .RESET_B(net1011),
    .SCD(net34),
    .SCE(net883),
    .Q(net858),
    .Q_N(net43));
 sky130_fd_sc_hd__a21bo_1 c111 (.A1(net788),
    .A2(net915),
    .B1_N(net818),
    .X(net867));
 sky130_fd_sc_hd__a21bo_1 c112 (.A1(net796),
    .A2(net3),
    .B1_N(net858),
    .X(net44));
 sky130_fd_sc_hd__buf_1 c113 (.A(net640),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 c114 (.A(net640),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 c115 (.A(net702),
    .X(net47));
 sky130_fd_sc_hd__xnor2_1 c116 (.A(net35),
    .B(net25),
    .Y(net48));
 sky130_fd_sc_hd__a21bo_1 c117 (.A1(net13),
    .A2(net47),
    .B1_N(net858),
    .X(net49));
 sky130_fd_sc_hd__xnor2_1 c118 (.A(net48),
    .B(net826),
    .Y(net50));
 sky130_fd_sc_hd__xnor2_1 c119 (.A(net4),
    .B(net883),
    .Y(net51));
 sky130_fd_sc_hd__xnor2_1 c120 (.A(net30),
    .B(net789),
    .Y(net52));
 sky130_fd_sc_hd__a41o_1 c121 (.A1(net50),
    .A2(net834),
    .A3(net800),
    .A4(net966),
    .B1(net15),
    .X(net53));
 sky130_fd_sc_hd__a31o_1 c122 (.A1(net51),
    .A2(net858),
    .A3(net799),
    .B1(net45),
    .X(net54));
 sky130_fd_sc_hd__xnor2_1 c123 (.A(net54),
    .B(net41),
    .Y(net880));
 sky130_fd_sc_hd__a41o_1 c124 (.A1(net53),
    .A2(net814),
    .A3(net966),
    .A4(net799),
    .B1(net34),
    .X(net55));
 sky130_fd_sc_hd__xnor2_2 c125 (.A(net45),
    .B(net809),
    .Y(net56));
 sky130_fd_sc_hd__xnor2_1 c126 (.A(net41),
    .B(net56),
    .Y(net57));
 sky130_fd_sc_hd__a21bo_2 c127 (.A1(net966),
    .A2(net880),
    .B1_N(net671),
    .X(net58));
 sky130_fd_sc_hd__a21bo_1 c128 (.A1(net15),
    .A2(net58),
    .B1_N(net41),
    .X(net59));
 sky130_fd_sc_hd__mux4_1 c129 (.A0(net46),
    .A1(net48),
    .A2(net58),
    .A3(net1001),
    .S0(net43),
    .S1(net56),
    .X(net60));
 sky130_fd_sc_hd__a21bo_1 c130 (.A1(net1009),
    .A2(net53),
    .B1_N(net58),
    .X(net891));
 sky130_fd_sc_hd__mux4_1 c131 (.A0(net59),
    .A1(net60),
    .A2(net891),
    .A3(net41),
    .S0(net58),
    .S1(net966),
    .X(net61));
 sky130_fd_sc_hd__xnor2_4 c132 (.A(net795),
    .B(net828),
    .Y(net62));
 sky130_fd_sc_hd__xnor2_4 c133 (.A(net644),
    .B(net817),
    .Y(net63));
 sky130_fd_sc_hd__xnor2_4 c134 (.A(net785),
    .B(net791),
    .Y(net64));
 sky130_fd_sc_hd__xnor2_4 c135 (.A(net63),
    .B(net1009),
    .Y(net65));
 sky130_fd_sc_hd__xnor2_4 c136 (.A(net999),
    .B(net930),
    .Y(net66));
 sky130_fd_sc_hd__xnor2_4 c137 (.A(net64),
    .B(net920),
    .Y(net67));
 sky130_fd_sc_hd__xnor2_4 c138 (.A(net960),
    .B(net794),
    .Y(net68));
 sky130_fd_sc_hd__xnor2_4 c139 (.A(net927),
    .B(net1006),
    .Y(net69));
 sky130_fd_sc_hd__xnor2_4 c140 (.A(net914),
    .B(net926),
    .Y(net70));
 sky130_fd_sc_hd__a21bo_4 c141 (.A1(net907),
    .A2(net926),
    .B1_N(net65),
    .X(net71));
 sky130_fd_sc_hd__xnor2_2 c142 (.A(net960),
    .B(net928),
    .Y(net72));
 sky130_fd_sc_hd__a21bo_4 c143 (.A1(net910),
    .A2(net920),
    .B1_N(net68),
    .X(net73));
 sky130_fd_sc_hd__a21bo_4 c144 (.A1(net928),
    .A2(net790),
    .B1_N(net909),
    .X(net74));
 sky130_fd_sc_hd__a41o_4 c145 (.A1(net905),
    .A2(net74),
    .A3(net66),
    .A4(net960),
    .B1(net909),
    .X(net75));
 sky130_fd_sc_hd__a21bo_4 c146 (.A1(net75),
    .A2(net806),
    .B1_N(net909),
    .X(net76));
 sky130_fd_sc_hd__xnor2_4 c147 (.A(net76),
    .B(net73),
    .Y(net77));
 sky130_fd_sc_hd__mux4_2 c148 (.A0(net69),
    .A1(net76),
    .A2(net77),
    .A3(net797),
    .S0(net785),
    .S1(net909),
    .X(net78));
 sky130_fd_sc_hd__a21bo_2 c149 (.A1(net905),
    .A2(net77),
    .B1_N(net907),
    .X(net79));
 sky130_fd_sc_hd__mux4_2 c150 (.A0(net806),
    .A1(net844),
    .A2(net909),
    .A3(net76),
    .S0(net960),
    .S1(net78),
    .X(net80));
 sky130_fd_sc_hd__a21bo_4 c151 (.A1(net902),
    .A2(net79),
    .B1_N(net909),
    .X(net81));
 sky130_fd_sc_hd__a41o_4 c152 (.A1(net902),
    .A2(net78),
    .A3(net77),
    .A4(net909),
    .B1(net74),
    .X(net82));
 sky130_fd_sc_hd__a21bo_4 c153 (.A1(net82),
    .A2(net992),
    .B1_N(net74),
    .X(net848));
 sky130_fd_sc_hd__xnor2_4 c154 (.A(net66),
    .B(net799),
    .Y(net83));
 sky130_fd_sc_hd__xnor2_4 c155 (.A(net798),
    .B(net67),
    .Y(net84));
 sky130_fd_sc_hd__xnor2_4 c156 (.A(net83),
    .B(net818),
    .Y(net85));
 sky130_fd_sc_hd__a21bo_4 c157 (.A1(net84),
    .A2(net811),
    .B1_N(net790),
    .X(net86));
 sky130_fd_sc_hd__a21bo_4 c158 (.A1(net816),
    .A2(net806),
    .B1_N(net799),
    .X(net87));
 sky130_fd_sc_hd__xnor2_4 c159 (.A(net800),
    .B(net908),
    .Y(net88));
 sky130_fd_sc_hd__a21bo_4 c160 (.A1(net809),
    .A2(net947),
    .B1_N(net86),
    .X(net89));
 sky130_fd_sc_hd__xnor2_4 c161 (.A(net87),
    .B(net790),
    .Y(net90));
 sky130_fd_sc_hd__xnor2_4 c162 (.A(net947),
    .B(net920),
    .Y(net857));
 sky130_fd_sc_hd__xnor2_4 c163 (.A(net90),
    .B(net813),
    .Y(net91));
 sky130_fd_sc_hd__xnor2_4 c164 (.A(net78),
    .B(net906),
    .Y(net92));
 sky130_fd_sc_hd__a21bo_2 c165 (.A1(net92),
    .A2(net818),
    .B1_N(net857),
    .X(net93));
 sky130_fd_sc_hd__mux4_2 c166 (.A0(net67),
    .A1(net90),
    .A2(net91),
    .A3(net88),
    .S0(net909),
    .S1(net83),
    .X(net94));
 sky130_fd_sc_hd__a21bo_4 c167 (.A1(net94),
    .A2(net92),
    .B1_N(net807),
    .X(net95));
 sky130_fd_sc_hd__xnor2_4 c168 (.A(net939),
    .B(net94),
    .Y(net96));
 sky130_fd_sc_hd__a21bo_4 c169 (.A1(net93),
    .A2(net96),
    .B1_N(net799),
    .X(net97));
 sky130_fd_sc_hd__a21bo_2 c170 (.A1(net92),
    .A2(net95),
    .B1_N(net88),
    .X(net98));
 sky130_fd_sc_hd__a31o_1 c171 (.A1(net98),
    .A2(net93),
    .A3(net97),
    .B1(net910),
    .X(net99));
 sky130_fd_sc_hd__mux4_2 c172 (.A0(net796),
    .A1(net91),
    .A2(net807),
    .A3(net1007),
    .S0(net906),
    .S1(net911),
    .X(net100));
 sky130_fd_sc_hd__xnor2_4 c173 (.A(net100),
    .B(net66),
    .Y(net101));
 sky130_fd_sc_hd__a21bo_2 c174 (.A1(net88),
    .A2(net790),
    .B1_N(net101),
    .X(net102));
 sky130_fd_sc_hd__mux4_2 c175 (.A0(net91),
    .A1(net94),
    .A2(net101),
    .A3(net82),
    .S0(net789),
    .S1(clknet_1_0__leaf_net693),
    .X(net103));
 sky130_fd_sc_hd__a21bo_2 c176 (.A1(net839),
    .A2(net93),
    .B1_N(net102),
    .X(net104));
 sky130_fd_sc_hd__xnor2_2 c177 (.A(net0),
    .B(net101),
    .Y(net105));
 sky130_fd_sc_hd__xnor2_2 c178 (.A(net929),
    .B(net906),
    .Y(net106));
 sky130_fd_sc_hd__buf_6 c179 (.A(clknet_1_1__leaf_net693),
    .X(net107));
 sky130_fd_sc_hd__a41o_2 c180 (.A1(net805),
    .A2(net806),
    .A3(net68),
    .A4(net809),
    .B1(net829),
    .X(net108));
 sky130_fd_sc_hd__a41o_2 c181 (.A1(net76),
    .A2(net108),
    .A3(net841),
    .A4(net84),
    .B1(net908),
    .X(net109));
 sky130_fd_sc_hd__a21bo_1 c182 (.A1(net101),
    .A2(net824),
    .B1_N(net911),
    .X(net110));
 sky130_fd_sc_hd__a21bo_1 c183 (.A1(net102),
    .A2(net68),
    .B1_N(net929),
    .X(net111));
 sky130_fd_sc_hd__a21bo_1 c184 (.A1(net96),
    .A2(net106),
    .B1_N(clknet_1_0__leaf_net693),
    .X(net112));
 sky130_fd_sc_hd__xnor2_4 c185 (.A(net830),
    .B(clknet_1_1__leaf_net107),
    .Y(net113));
 sky130_fd_sc_hd__a21bo_1 c186 (.A1(clknet_1_0__leaf_net112),
    .A2(net111),
    .B1_N(net825),
    .X(net114));
 sky130_fd_sc_hd__xnor2_1 c187 (.A(net108),
    .B(net79),
    .Y(net115));
 sky130_fd_sc_hd__a21bo_1 c188 (.A1(net0),
    .A2(net911),
    .B1_N(clknet_1_1__leaf_net693),
    .X(net116));
 sky130_fd_sc_hd__buf_1 c189 (.A(clknet_1_0__leaf_net693),
    .X(net117));
 sky130_fd_sc_hd__a21bo_1 c190 (.A1(clknet_1_0__leaf_net107),
    .A2(clknet_1_0__leaf_net117),
    .B1_N(clknet_1_0__leaf_net113),
    .X(net118));
 sky130_fd_sc_hd__xnor2_1 c191 (.A(clknet_1_1__leaf_net113),
    .B(net115),
    .Y(net119));
 sky130_fd_sc_hd__mux4_2 c192 (.A0(clknet_1_0__leaf_net118),
    .A1(net95),
    .A2(net1010),
    .A3(net86),
    .S0(net835),
    .S1(net110),
    .X(net120));
 sky130_fd_sc_hd__buf_1 c193 (.A(clknet_1_1__leaf_net693),
    .X(net121));
 sky130_fd_sc_hd__a21bo_1 c194 (.A1(clknet_1_0__leaf_net120),
    .A2(net100),
    .B1_N(clknet_1_1__leaf_net119),
    .X(net122));
 sky130_fd_sc_hd__a31o_1 c195 (.A1(net111),
    .A2(net73),
    .A3(net829),
    .B1(net89),
    .X(net123));
 sky130_fd_sc_hd__mux4_1 c196 (.A0(net106),
    .A1(net108),
    .A2(clknet_1_0__leaf_net117),
    .A3(net841),
    .S0(net123),
    .S1(clknet_1_0__leaf_net118),
    .X(net124));
 sky130_fd_sc_hd__a21bo_1 c197 (.A1(clknet_1_0__leaf_net122),
    .A2(net68),
    .B1_N(net123),
    .X(net125));
 sky130_fd_sc_hd__a21bo_1 c198 (.A1(net18),
    .A2(clknet_1_1__leaf_net119),
    .B1_N(net791),
    .X(net126));
 sky130_fd_sc_hd__a21bo_1 c199 (.A1(net795),
    .A2(net829),
    .B1_N(clknet_1_0__leaf_net122),
    .X(net127));
 sky130_fd_sc_hd__buf_2 c200 (.A(net887),
    .X(net128));
 sky130_fd_sc_hd__a31o_4 c201 (.A1(clknet_1_1__leaf_net118),
    .A2(net791),
    .A3(net17),
    .B1(net917),
    .X(net129));
 sky130_fd_sc_hd__a21bo_1 c202 (.A1(net94),
    .A2(net2),
    .B1_N(net926),
    .X(net130));
 sky130_fd_sc_hd__buf_1 c203 (.A(net887),
    .X(net131));
 sky130_fd_sc_hd__a21bo_1 c204 (.A1(clknet_1_1__leaf_net118),
    .A2(net805),
    .B1_N(net130),
    .X(net132));
 sky130_fd_sc_hd__mux4_1 c205 (.A0(clknet_1_0__leaf_net129),
    .A1(clknet_1_0__leaf_net127),
    .A2(net14),
    .A3(net9),
    .S0(net798),
    .S1(net917),
    .X(net133));
 sky130_fd_sc_hd__a41o_1 c206 (.A1(clknet_1_1__leaf_net129),
    .A2(net17),
    .A3(net18),
    .A4(clknet_1_0__leaf_net132),
    .B1(net917),
    .X(net134));
 sky130_fd_sc_hd__mux4_2 c207 (.A0(net930),
    .A1(net105),
    .A2(net928),
    .A3(net916),
    .S0(net3),
    .S1(net795),
    .X(net135));
 sky130_fd_sc_hd__a41o_1 c208 (.A1(net11),
    .A2(net135),
    .A3(clknet_1_0__leaf_net126),
    .A4(net918),
    .B1(net916),
    .X(net136));
 sky130_fd_sc_hd__a21bo_1 c209 (.A1(clknet_1_0__leaf_net134),
    .A2(net2),
    .B1_N(net976),
    .X(net137));
 sky130_fd_sc_hd__mux4_1 c210 (.A0(net824),
    .A1(clknet_1_0__leaf_net127),
    .A2(clknet_1_0__leaf_net129),
    .A3(clknet_1_0__leaf_net119),
    .S0(net820),
    .S1(net917),
    .X(net138));
 sky130_fd_sc_hd__mux4_1 c211 (.A0(clknet_1_0__leaf_net119),
    .A1(net3),
    .A2(net98),
    .A3(clknet_1_0__leaf_net136),
    .S0(clknet_1_0__leaf_net129),
    .S1(net917),
    .X(net139));
 sky130_fd_sc_hd__a21bo_1 c212 (.A1(net111),
    .A2(clknet_1_0__leaf_net132),
    .B1_N(clknet_1_0__leaf_net134),
    .X(net140));
 sky130_fd_sc_hd__a21bo_2 c213 (.A1(net9),
    .A2(net805),
    .B1_N(net799),
    .X(net141));
 sky130_fd_sc_hd__a41o_1 c214 (.A1(clknet_1_0__leaf_net134),
    .A2(net839),
    .A3(clknet_1_0__leaf_net140),
    .A4(net917),
    .B1(net79),
    .X(net142));
 sky130_fd_sc_hd__a41o_1 c215 (.A1(clknet_1_0__leaf_net142),
    .A2(net18),
    .A3(net796),
    .A4(clknet_1_0__leaf_net134),
    .B1(clknet_1_0__leaf_net140),
    .X(net143));
 sky130_fd_sc_hd__mux4_1 c216 (.A0(net115),
    .A1(net79),
    .A2(clknet_1_1__leaf_net136),
    .A3(clknet_1_0__leaf_net137),
    .S0(clknet_1_0__leaf_net140),
    .S1(net815),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 c217 (.A(net702),
    .X(net876));
 sky130_fd_sc_hd__sdfbbn_1 c218 (.CLK_N(clknet_4_1_0_clk),
    .D(clknet_1_0__leaf_net144),
    .RESET_B(clknet_1_0__leaf_net143),
    .SCD(net21),
    .SCE(clknet_1_0__leaf_net134),
    .SET_B(net917),
    .Q(net146),
    .Q_N(net145));
 sky130_fd_sc_hd__sdfrtn_1 c219 (.CLK_N(clknet_4_1_0_clk),
    .D(net917),
    .RESET_B(net21),
    .SCD(clknet_1_1__leaf_net144),
    .SCE(net911),
    .Q(net147));
 sky130_fd_sc_hd__a21bo_1 c220 (.A1(net835),
    .A2(net908),
    .B1_N(net806),
    .X(net148));
 sky130_fd_sc_hd__a21bo_1 c221 (.A1(net14),
    .A2(net33),
    .B1_N(clknet_1_0__leaf_net142),
    .X(net149));
 sky130_fd_sc_hd__a21bo_1 c222 (.A1(net10),
    .A2(net922),
    .B1_N(net6),
    .X(net150));
 sky130_fd_sc_hd__sdfrtp_2 c223 (.CLK(clknet_4_4_0_clk),
    .D(net105),
    .RESET_B(clknet_1_0__leaf_net149),
    .SCD(clknet_1_0__leaf_net126),
    .SCE(clknet_1_1__leaf_net693),
    .Q(net151));
 sky130_fd_sc_hd__a21bo_1 c224 (.A1(net25),
    .A2(net810),
    .B1_N(net922),
    .X(net152));
 sky130_fd_sc_hd__buf_1 c225 (.A(net703),
    .X(net153));
 sky130_fd_sc_hd__a31o_1 c226 (.A1(net105),
    .A2(clknet_1_0__leaf_net139),
    .A3(net89),
    .B1(net930),
    .X(net154));
 sky130_fd_sc_hd__a21bo_1 c227 (.A1(net38),
    .A2(net976),
    .B1_N(net675),
    .X(net155));
 sky130_fd_sc_hd__a21bo_1 c228 (.A1(net29),
    .A2(net153),
    .B1_N(net148),
    .X(net156));
 sky130_fd_sc_hd__a21bo_2 c229 (.A1(net794),
    .A2(net81),
    .B1_N(net27),
    .X(net157));
 sky130_fd_sc_hd__a31o_2 c230 (.A1(net95),
    .A2(net157),
    .A3(net857),
    .B1(net28),
    .X(net158));
 sky130_fd_sc_hd__a21bo_2 c231 (.A1(net821),
    .A2(net105),
    .B1_N(net158),
    .X(net159));
 sky130_fd_sc_hd__a31o_2 c232 (.A1(net155),
    .A2(net135),
    .A3(net150),
    .B1(net158),
    .X(net856));
 sky130_fd_sc_hd__a41o_1 c233 (.A1(clknet_1_1__leaf_net129),
    .A2(net807),
    .A3(net153),
    .A4(net158),
    .B1(net896),
    .X(net160));
 sky130_fd_sc_hd__mux4_2 c234 (.A0(net12),
    .A1(net821),
    .A2(net834),
    .A3(net922),
    .S0(net980),
    .S1(net911),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 c235 (.A(net703),
    .X(net162));
 sky130_fd_sc_hd__sdfrtp_1 c236 (.CLK(clknet_4_4_0_clk),
    .D(net156),
    .RESET_B(net109),
    .SCD(net158),
    .SCE(net896),
    .Q(net163));
 sky130_fd_sc_hd__mux4_1 c237 (.A0(net976),
    .A1(net159),
    .A2(net896),
    .A3(net155),
    .S0(net141),
    .S1(net675),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_2 c238 (.A(net702),
    .X(net851));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(clknet_1_1__leaf_net139),
    .A1(net158),
    .A2(net162),
    .A3(net896),
    .S0(net163),
    .S1(net155),
    .X(net165));
 sky130_fd_sc_hd__a31o_1 c240 (.A1(net157),
    .A2(net162),
    .A3(net918),
    .B1(net701),
    .X(net166));
 sky130_fd_sc_hd__a41o_1 c241 (.A1(net153),
    .A2(net163),
    .A3(net166),
    .A4(net896),
    .X(net167));
 sky130_fd_sc_hd__a21bo_1 c242 (.A1(net3),
    .A2(net834),
    .B1_N(net671),
    .X(net168));
 sky130_fd_sc_hd__a31o_1 c243 (.A1(net28),
    .A2(net58),
    .A3(net896),
    .B1(net795),
    .X(net169));
 sky130_fd_sc_hd__a21bo_1 c244 (.A1(net93),
    .A2(net109),
    .B1_N(clknet_1_1__leaf_net126),
    .X(net170));
 sky130_fd_sc_hd__a21bo_1 c245 (.A1(net52),
    .A2(net168),
    .B1_N(net867),
    .X(net888));
 sky130_fd_sc_hd__a31o_1 c246 (.A1(net44),
    .A2(net109),
    .A3(clknet_1_1__leaf_net170),
    .B1(net58),
    .X(net171));
 sky130_fd_sc_hd__a41o_1 c247 (.A1(net834),
    .A2(net49),
    .A3(net888),
    .A4(net883),
    .B1(net671),
    .X(net172));
 sky130_fd_sc_hd__a31o_1 c248 (.A1(clknet_1_1__leaf_net126),
    .A2(net28),
    .A3(net52),
    .B1(net56),
    .X(net884));
 sky130_fd_sc_hd__a31o_1 c249 (.A1(net47),
    .A2(net796),
    .A3(net44),
    .B1(net43),
    .X(net889));
 sky130_fd_sc_hd__mux4_1 c250 (.A0(clknet_1_0__leaf_net170),
    .A1(clknet_1_0__leaf_net884),
    .A2(net860),
    .A3(net58),
    .S0(net915),
    .S1(net710),
    .X(net173));
 sky130_fd_sc_hd__a21bo_1 c251 (.A1(net3),
    .A2(net848),
    .B1_N(net712),
    .X(net174));
 sky130_fd_sc_hd__a41o_1 c252 (.A1(net800),
    .A2(clknet_1_1__leaf_net884),
    .A3(net881),
    .A4(net709),
    .B1(net712),
    .X(net175));
 sky130_fd_sc_hd__a21bo_1 c253 (.A1(net109),
    .A2(net872),
    .B1_N(net883),
    .X(net176));
 sky130_fd_sc_hd__mux4_1 c254 (.A0(net172),
    .A1(net915),
    .A2(net176),
    .A3(net90),
    .S0(clknet_1_1__leaf_net884),
    .S1(net712),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 c255 (.A0(net807),
    .A1(net47),
    .A2(net176),
    .A3(net25),
    .S0(net671),
    .S1(net710),
    .X(net178));
 sky130_fd_sc_hd__a21bo_1 c256 (.A1(net178),
    .A2(net176),
    .B1_N(net860),
    .X(net865));
 sky130_fd_sc_hd__a21bo_1 c257 (.A1(net90),
    .A2(net176),
    .B1_N(net858),
    .X(net179));
 sky130_fd_sc_hd__buf_1 c258 (.A(net781),
    .X(net861));
 sky130_fd_sc_hd__sdfbbn_1 c259 (.CLK_N(clknet_4_5_0_clk),
    .D(net174),
    .RESET_B(net56),
    .SCD(clknet_1_1__leaf_net126),
    .SCE(net896),
    .SET_B(net865),
    .Q(net885),
    .Q_N(net180));
 sky130_fd_sc_hd__mux4_1 c260 (.A0(net97),
    .A1(net179),
    .A2(net58),
    .A3(net915),
    .S0(net43),
    .S1(net25),
    .X(net181));
 sky130_fd_sc_hd__a21bo_1 c261 (.A1(net846),
    .A2(net889),
    .B1_N(net710),
    .X(net182));
 sky130_fd_sc_hd__mux4_1 c262 (.A0(net176),
    .A1(net785),
    .A2(net182),
    .A3(net180),
    .S0(net881),
    .S1(net711),
    .X(net183));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net183),
    .A1(net182),
    .A2(net861),
    .A3(net56),
    .S0(net709),
    .S1(net711),
    .X(net184));
 sky130_fd_sc_hd__a21bo_4 c264 (.A1(net794),
    .A2(net839),
    .B1_N(net77),
    .X(net185));
 sky130_fd_sc_hd__xnor2_4 c265 (.A(net791),
    .B(net954),
    .Y(net186));
 sky130_fd_sc_hd__xnor2_4 c266 (.A(net186),
    .B(net951),
    .Y(net187));
 sky130_fd_sc_hd__xnor2_4 c267 (.A(net795),
    .B(net913),
    .Y(net188));
 sky130_fd_sc_hd__a21bo_2 c268 (.A1(net790),
    .A2(net828),
    .B1_N(net81),
    .X(net189));
 sky130_fd_sc_hd__xnor2_4 c269 (.A(net185),
    .B(net934),
    .Y(net190));
 sky130_fd_sc_hd__xnor2_2 c270 (.A(net188),
    .B(net187),
    .Y(net191));
 sky130_fd_sc_hd__xnor2_4 c271 (.A(net913),
    .B(net70),
    .Y(net192));
 sky130_fd_sc_hd__xnor2_4 c272 (.A(net935),
    .B(net900),
    .Y(net193));
 sky130_fd_sc_hd__xnor2_4 c273 (.A(net192),
    .B(net188),
    .Y(net194));
 sky130_fd_sc_hd__xnor2_4 c274 (.A(net900),
    .B(net193),
    .Y(net195));
 sky130_fd_sc_hd__xnor2_1 c275 (.A(net187),
    .B(net898),
    .Y(net196));
 sky130_fd_sc_hd__a21bo_4 c276 (.A1(net190),
    .A2(net902),
    .B1_N(net900),
    .X(net197));
 sky130_fd_sc_hd__xnor2_4 c277 (.A(net197),
    .B(net903),
    .Y(net198));
 sky130_fd_sc_hd__xnor2_4 c278 (.A(net898),
    .B(net198),
    .Y(net853));
 sky130_fd_sc_hd__clkbuf_2 c279 (.A(net707),
    .X(net199));
 sky130_fd_sc_hd__a21bo_4 c280 (.A1(net189),
    .A2(net190),
    .B1_N(net828),
    .X(net200));
 sky130_fd_sc_hd__a21bo_4 c281 (.A1(net194),
    .A2(net187),
    .B1_N(net199),
    .X(net201));
 sky130_fd_sc_hd__a21bo_1 c282 (.A1(net201),
    .A2(net790),
    .B1_N(net198),
    .X(net202));
 sky130_fd_sc_hd__a21bo_2 c283 (.A1(net200),
    .A2(net192),
    .B1_N(net74),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_8 c284 (.A(net707),
    .X(net870));
 sky130_fd_sc_hd__a21bo_1 c285 (.A1(net74),
    .A2(net870),
    .B1_N(net188),
    .X(net204));
 sky130_fd_sc_hd__xnor2_4 c286 (.A(net190),
    .B(net88),
    .Y(net205));
 sky130_fd_sc_hd__xnor2_2 c287 (.A(net86),
    .B(net931),
    .Y(net206));
 sky130_fd_sc_hd__a21bo_2 c288 (.A1(net931),
    .A2(net205),
    .B1_N(net907),
    .X(net207));
 sky130_fd_sc_hd__xnor2_4 c289 (.A(net815),
    .B(net816),
    .Y(net877));
 sky130_fd_sc_hd__a31o_2 c290 (.A1(net66),
    .A2(net199),
    .A3(net87),
    .B1(net909),
    .X(net208));
 sky130_fd_sc_hd__xnor2_4 c291 (.A(net186),
    .B(net870),
    .Y(net209));
 sky130_fd_sc_hd__a21bo_4 c292 (.A1(net208),
    .A2(net804),
    .B1_N(net813),
    .X(net210));
 sky130_fd_sc_hd__xnor2_2 c293 (.A(net857),
    .B(net88),
    .Y(net874));
 sky130_fd_sc_hd__xnor2_4 c294 (.A(net897),
    .B(net870),
    .Y(net211));
 sky130_fd_sc_hd__a31o_1 c295 (.A1(net211),
    .A2(net102),
    .A3(net794),
    .B1(net83),
    .X(net212));
 sky130_fd_sc_hd__xnor2_4 c296 (.A(net804),
    .B(net925),
    .Y(net213));
 sky130_fd_sc_hd__xnor2_2 c297 (.A(net205),
    .B(net208),
    .Y(net214));
 sky130_fd_sc_hd__a21bo_4 c298 (.A1(net214),
    .A2(net815),
    .B1_N(net210),
    .X(net215));
 sky130_fd_sc_hd__mux4_1 c299 (.A0(net209),
    .A1(net211),
    .A2(net185),
    .A3(net820),
    .S0(net926),
    .S1(net877),
    .X(net216));
 sky130_fd_sc_hd__xnor2_4 c300 (.A(net86),
    .B(net804),
    .Y(net217));
 sky130_fd_sc_hd__a41o_1 c301 (.A1(net217),
    .A2(net186),
    .A3(net78),
    .A4(net692),
    .B1(net713),
    .X(net218));
 sky130_fd_sc_hd__xnor2_4 c302 (.A(net215),
    .B(net206),
    .Y(net219));
 sky130_fd_sc_hd__xnor2_1 c303 (.A(net814),
    .B(net205),
    .Y(net220));
 sky130_fd_sc_hd__mux4_1 c304 (.A0(net218),
    .A1(net219),
    .A2(net220),
    .A3(net900),
    .S0(net84),
    .S1(net211),
    .X(net221));
 sky130_fd_sc_hd__a41o_1 c305 (.A1(net199),
    .A2(net217),
    .A3(net909),
    .A4(net691),
    .B1(net713),
    .X(net222));
 sky130_fd_sc_hd__a21bo_1 c306 (.A1(net88),
    .A2(net222),
    .B1_N(net691),
    .X(net223));
 sky130_fd_sc_hd__mux4_2 c307 (.A0(net204),
    .A1(net220),
    .A2(net223),
    .A3(net66),
    .S0(net199),
    .S1(net691),
    .X(net224));
 sky130_fd_sc_hd__a31o_1 c308 (.A1(clknet_1_0__leaf_net125),
    .A2(clknet_1_1__leaf_net112),
    .A3(clknet_1_0__leaf_net122),
    .B1(net897),
    .X(net225));
 sky130_fd_sc_hd__a31o_1 c309 (.A1(net930),
    .A2(net86),
    .A3(net825),
    .B1(clknet_1_1__leaf_net114),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_2 c310 (.A(net776),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_4 c311 (.A(net776),
    .X(net228));
 sky130_fd_sc_hd__mux4_1 c312 (.A0(net934),
    .A1(net877),
    .A2(net853),
    .A3(clknet_1_0__leaf_net112),
    .S0(net185),
    .S1(net819),
    .X(net229));
 sky130_fd_sc_hd__xnor2_1 c313 (.A(clknet_1_0__leaf_net107),
    .B(clknet_1_0__leaf_net121),
    .Y(net230));
 sky130_fd_sc_hd__xnor2_2 c314 (.A(net98),
    .B(net979),
    .Y(net231));
 sky130_fd_sc_hd__mux4_2 c315 (.A0(net940),
    .A1(clknet_1_1__leaf_net117),
    .A2(clknet_1_1__leaf_net230),
    .A3(clknet_1_0__leaf_net120),
    .S0(net228),
    .S1(net110),
    .X(net232));
 sky130_fd_sc_hd__xnor2_4 c316 (.A(net811),
    .B(clknet_1_0__leaf_net232),
    .Y(net233));
 sky130_fd_sc_hd__a21bo_2 c317 (.A1(net106),
    .A2(net210),
    .B1_N(net123),
    .X(net234));
 sky130_fd_sc_hd__xnor2_1 c318 (.A(net110),
    .B(net231),
    .Y(net235));
 sky130_fd_sc_hd__a21bo_2 c319 (.A1(net220),
    .A2(net897),
    .B1_N(net910),
    .X(net236));
 sky130_fd_sc_hd__buf_1 c320 (.A(clknet_1_0__leaf_net693),
    .X(net237));
 sky130_fd_sc_hd__a21bo_1 c321 (.A1(net187),
    .A2(net832),
    .B1_N(net691),
    .X(net238));
 sky130_fd_sc_hd__a21bo_1 c322 (.A1(clknet_1_0__leaf_net113),
    .A2(net223),
    .B1_N(net910),
    .X(net239));
 sky130_fd_sc_hd__mux4_1 c323 (.A0(clknet_1_0__leaf_net233),
    .A1(net897),
    .A2(net841),
    .A3(net189),
    .S0(net236),
    .S1(net234),
    .X(net240));
 sky130_fd_sc_hd__buf_2 c324 (.A(net778),
    .X(net869));
 sky130_fd_sc_hd__a21bo_1 c325 (.A1(clknet_1_0__leaf_net237),
    .A2(clknet_1_0__leaf_net122),
    .B1_N(net840),
    .X(net241));
 sky130_fd_sc_hd__buf_1 c326 (.A(net690),
    .X(net242));
 sky130_fd_sc_hd__xnor2_2 c327 (.A(net842),
    .B(net210),
    .Y(net243));
 sky130_fd_sc_hd__dfbbn_1 c328 (.CLK_N(clknet_4_2_0_clk),
    .D(clknet_1_0__leaf_net241),
    .RESET_B(net231),
    .SET_B(net243),
    .Q(net245),
    .Q_N(net244));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net245),
    .A1(clknet_1_1__leaf_net241),
    .A2(net243),
    .A3(clknet_1_0__leaf_net239),
    .S0(net234),
    .S1(net201),
    .X(net246));
 sky130_fd_sc_hd__a31o_1 c330 (.A1(net244),
    .A2(net8),
    .A3(net193),
    .B1(net832),
    .X(net247));
 sky130_fd_sc_hd__a31o_1 c331 (.A1(net247),
    .A2(net823),
    .A3(net200),
    .B1(net930),
    .X(net248));
 sky130_fd_sc_hd__a41o_1 c332 (.A1(net925),
    .A2(net228),
    .A3(net69),
    .A4(net839),
    .B1(clknet_1_0__leaf_net716),
    .X(net249));
 sky130_fd_sc_hd__a31o_1 c333 (.A1(net243),
    .A2(clknet_1_1__leaf_net249),
    .A3(net1004),
    .B1(net185),
    .X(net250));
 sky130_fd_sc_hd__a21bo_1 c334 (.A1(clknet_1_0__leaf_net112),
    .A2(net818),
    .B1_N(clknet_1_0__leaf_net715),
    .X(net251));
 sky130_fd_sc_hd__a21bo_1 c335 (.A1(net208),
    .A2(net79),
    .B1_N(net247),
    .X(net252));
 sky130_fd_sc_hd__sdfbbp_1 c336 (.CLK(clknet_4_0_0_clk),
    .D(clknet_1_0__leaf_net249),
    .RESET_B(clknet_1_0__leaf_net127),
    .SCD(net877),
    .SCE(net17),
    .SET_B(net887),
    .Q(net254),
    .Q_N(net253));
 sky130_fd_sc_hd__sdfrtp_1 c337 (.CLK(clknet_4_1_0_clk),
    .D(clknet_1_1__leaf_net143),
    .RESET_B(clknet_1_0__leaf_net251),
    .SCD(clknet_1_1__leaf_net137),
    .SCE(net898),
    .Q(net255));
 sky130_fd_sc_hd__a31o_1 c338 (.A1(net254),
    .A2(net959),
    .A3(clknet_1_0__leaf_net233),
    .B1(net703),
    .X(net256));
 sky130_fd_sc_hd__a31o_1 c339 (.A1(net234),
    .A2(net84),
    .A3(net897),
    .B1(net905),
    .X(net257));
 sky130_fd_sc_hd__a41o_1 c340 (.A1(net84),
    .A2(net63),
    .A3(net253),
    .A4(net108),
    .B1(net860),
    .X(net258));
 sky130_fd_sc_hd__sdfsbp_1 c341 (.CLK(clknet_4_0_0_clk),
    .D(clknet_1_0__leaf_net251),
    .SCD(clknet_1_0__leaf_net136),
    .SCE(net667),
    .SET_B(clknet_1_1__leaf_net715),
    .Q(net260),
    .Q_N(net259));
 sky130_fd_sc_hd__clkbuf_1 c342 (.X(net261));
 sky130_fd_sc_hd__buf_1 c343 (.A(net643),
    .X(net892));
 sky130_fd_sc_hd__clkbuf_1 c344 (.A(net702),
    .X(net262));
 sky130_fd_sc_hd__a21bo_1 c345 (.A1(net892),
    .A2(clknet_1_0__leaf_net137),
    .B1_N(net141),
    .X(net263));
 sky130_fd_sc_hd__sdfbbn_1 c346 (.CLK_N(clknet_4_1_0_clk),
    .D(net9),
    .RESET_B(net876),
    .SCD(clknet_1_0__leaf_net251),
    .SCE(clknet_1_1__leaf_net249),
    .SET_B(net979),
    .Q(net265),
    .Q_N(net264));
 sky130_fd_sc_hd__a41o_1 c347 (.A1(net79),
    .A2(net261),
    .A3(clknet_1_1__leaf_net249),
    .A4(net832),
    .B1(net243),
    .X(net266));
 sky130_fd_sc_hd__mux4_1 c348 (.A0(net260),
    .A1(clknet_1_0__leaf_net121),
    .A2(clknet_1_0__leaf_net249),
    .A3(net252),
    .S0(net6),
    .S1(net236),
    .X(net267));
 sky130_fd_sc_hd__a41o_4 c349 (.A1(clknet_1_0__leaf_net263),
    .A2(net265),
    .A3(net147),
    .A4(net829),
    .B1(net259),
    .X(net268));
 sky130_fd_sc_hd__a41o_1 c350 (.A1(net198),
    .A2(clknet_1_0__leaf_net266),
    .A3(net264),
    .A4(net952),
    .B1(net886),
    .X(net269));
 sky130_fd_sc_hd__a31o_1 c351 (.A1(clknet_1_1__leaf_net266),
    .A2(clknet_1_0__leaf_net268),
    .A3(net258),
    .B1(clknet_1_1__leaf_net263),
    .X(net270));
 sky130_fd_sc_hd__sdfbbn_1 c352 (.CLK_N(clknet_4_4_0_clk),
    .D(net130),
    .RESET_B(net141),
    .SCD(net97),
    .SCE(net152),
    .SET_B(net701),
    .Q(net272),
    .Q_N(net271));
 sky130_fd_sc_hd__mux4_1 c353 (.A0(net150),
    .A1(net32),
    .A2(net876),
    .A3(net238),
    .S0(net922),
    .S1(net911),
    .X(net273));
 sky130_fd_sc_hd__a41o_1 c354 (.A1(net98),
    .A2(net79),
    .A3(net995),
    .A4(net813),
    .B1(net870),
    .X(net274));
 sky130_fd_sc_hd__a41o_2 c355 (.A1(net16),
    .A2(net101),
    .A3(net209),
    .A4(net271),
    .B1(net274),
    .X(net275));
 sky130_fd_sc_hd__a41o_2 c356 (.A1(net130),
    .A2(net918),
    .A3(net876),
    .A4(net995),
    .B1(net161),
    .X(net276));
 sky130_fd_sc_hd__a41o_2 c357 (.A1(net258),
    .A2(net148),
    .A3(net975),
    .A4(net38),
    .B1(net904),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 c358 (.A0(net162),
    .A1(net92),
    .A2(net928),
    .A3(net786),
    .S0(net911),
    .S1(net701),
    .X(net278));
 sky130_fd_sc_hd__a41o_1 c359 (.A1(clknet_1_1__leaf_net121),
    .A2(clknet_1_1__leaf_net230),
    .A3(net272),
    .A4(net219),
    .B1(net803),
    .X(net279));
 sky130_fd_sc_hd__a41o_1 c360 (.A1(net273),
    .A2(net157),
    .A3(net1003),
    .A4(net832),
    .B1(net688),
    .X(net280));
 sky130_fd_sc_hd__mux4_1 c361 (.A0(net815),
    .A1(net102),
    .A2(net258),
    .A3(net277),
    .S0(net932),
    .S1(net911),
    .X(net281));
 sky130_fd_sc_hd__a41o_1 c362 (.A1(net238),
    .A2(net272),
    .A3(net146),
    .A4(net846),
    .B1(clknet_1_0__leaf_net142),
    .X(net282));
 sky130_fd_sc_hd__sdfbbp_1 c363 (.CLK(clknet_4_6_0_clk),
    .D(net281),
    .RESET_B(net162),
    .SCD(net897),
    .SCE(net952),
    .SET_B(net275),
    .Q(net284),
    .Q_N(net283));
 sky130_fd_sc_hd__a41o_1 c364 (.A1(net975),
    .A2(net852),
    .A3(net275),
    .A4(net908),
    .B1(net281),
    .X(net285));
 sky130_fd_sc_hd__mux4_1 c365 (.A0(net788),
    .A1(net837),
    .A2(net278),
    .A3(clknet_1_1__leaf_net230),
    .S0(net161),
    .S1(net896),
    .X(net286));
 sky130_fd_sc_hd__sdfbbn_1 c366 (.CLK_N(clknet_4_4_0_clk),
    .D(net883),
    .RESET_B(clknet_1_1__leaf_net251),
    .SCD(net101),
    .SCE(net277),
    .SET_B(net688),
    .Q(net288),
    .Q_N(net287));
 sky130_fd_sc_hd__a41o_1 c367 (.A1(net280),
    .A2(net193),
    .A3(clknet_1_1__leaf_net134),
    .A4(net287),
    .B1(clknet_1_0__leaf_net863),
    .X(net289));
 sky130_fd_sc_hd__a41o_1 c368 (.A1(net817),
    .A2(net150),
    .A3(net157),
    .A4(net922),
    .B1(clknet_1_0__leaf_net863),
    .X(net290));
 sky130_fd_sc_hd__a41o_1 c369 (.A1(net278),
    .A2(net277),
    .A3(net813),
    .A4(net883),
    .B1(clknet_1_0__leaf_net863),
    .X(net291));
 sky130_fd_sc_hd__mux4_1 c370 (.A0(net274),
    .A1(net291),
    .A2(net843),
    .A3(clknet_1_0__leaf_net290),
    .S0(net1003),
    .S1(clknet_1_1__leaf_net863),
    .X(net292));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(net91),
    .A1(net275),
    .A2(net843),
    .A3(net283),
    .S0(clknet_1_0__leaf_net292),
    .S1(clknet_1_0__leaf_net863),
    .X(net293));
 sky130_fd_sc_hd__a41o_1 c372 (.A1(net163),
    .A2(net162),
    .A3(net869),
    .A4(net38),
    .B1(net717),
    .X(net882));
 sky130_fd_sc_hd__sdfbbn_2 c373 (.CLK_N(clknet_4_5_0_clk),
    .D(net6),
    .RESET_B(net289),
    .SCD(net872),
    .SCE(clknet_1_0__leaf_net292),
    .SET_B(clknet_1_1__leaf_net134),
    .Q(net295),
    .Q_N(net294));
 sky130_fd_sc_hd__mux4_1 c392 (.A0(net189),
    .A1(net177),
    .A2(net97),
    .A3(net814),
    .S0(net846),
    .S1(net882),
    .X(net296));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net168),
    .A1(clknet_1_0__leaf_net269),
    .A2(net184),
    .A3(clknet_1_1__leaf_net292),
    .S0(net856),
    .S1(net859),
    .X(net297));
 sky130_fd_sc_hd__mux4_1 c394 (.A0(net58),
    .A1(clknet_1_1__leaf_net292),
    .A2(net846),
    .A3(clknet_1_1__leaf_net269),
    .S0(net925),
    .S1(net719),
    .X(net298));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net800),
    .A1(net57),
    .A2(net58),
    .A3(clknet_1_0__leaf_net269),
    .S0(net851),
    .S1(net848),
    .X(net299));
 sky130_fd_sc_hd__buf_2 c396 (.A(net669),
    .X(net300));
 sky130_fd_sc_hd__buf_4 c397 (.A(net669),
    .X(net301));
 sky130_fd_sc_hd__xnor2_4 c398 (.A(net997),
    .B(net301),
    .Y(net302));
 sky130_fd_sc_hd__clkbuf_4 c399 (.A(net986),
    .X(net303));
 sky130_fd_sc_hd__xnor2_4 c400 (.A(net903),
    .B(net303),
    .Y(net849));
 sky130_fd_sc_hd__xnor2_1 c401 (.A(net192),
    .B(net198),
    .Y(net304));
 sky130_fd_sc_hd__xnor2_4 c402 (.A(net644),
    .B(net201),
    .Y(net305));
 sky130_fd_sc_hd__a21bo_4 c403 (.A1(net204),
    .A2(net301),
    .B1_N(net903),
    .X(net306));
 sky130_fd_sc_hd__xnor2_2 c404 (.A(net305),
    .B(net301),
    .Y(net307));
 sky130_fd_sc_hd__xnor2_2 c405 (.A(net300),
    .B(net74),
    .Y(net871));
 sky130_fd_sc_hd__xnor2_4 c406 (.A(net306),
    .B(net839),
    .Y(net308));
 sky130_fd_sc_hd__xnor2_2 c407 (.A(net307),
    .B(net302),
    .Y(net309));
 sky130_fd_sc_hd__a21bo_1 c408 (.A1(net955),
    .A2(net303),
    .B1_N(net910),
    .X(net310));
 sky130_fd_sc_hd__a21bo_1 c409 (.A1(net849),
    .A2(net956),
    .B1_N(net905),
    .X(net311));
 sky130_fd_sc_hd__xnor2_4 c410 (.A(net308),
    .B(net306),
    .Y(net312));
 sky130_fd_sc_hd__buf_1 c411 (.A(net778),
    .X(net313));
 sky130_fd_sc_hd__a21bo_1 c412 (.A1(net871),
    .A2(net307),
    .B1_N(net786),
    .X(net314));
 sky130_fd_sc_hd__a21bo_2 c413 (.A1(net310),
    .A2(net313),
    .B1_N(net905),
    .X(net315));
 sky130_fd_sc_hd__a41o_1 c414 (.A1(net313),
    .A2(net309),
    .A3(net849),
    .A4(net871),
    .B1(net305),
    .X(net316));
 sky130_fd_sc_hd__a21bo_4 c415 (.A1(net303),
    .A2(net315),
    .B1_N(net669),
    .X(net317));
 sky130_fd_sc_hd__a21bo_2 c416 (.A1(net315),
    .A2(net317),
    .B1_N(net910),
    .X(net318));
 sky130_fd_sc_hd__sdfbbp_1 c417 (.CLK(clknet_4_8_0_clk),
    .D(net314),
    .RESET_B(net204),
    .SCD(net303),
    .SCE(net317),
    .SET_B(net310),
    .Q(net320),
    .Q_N(net319));
 sky130_fd_sc_hd__clkbuf_2 c418 (.A(net690),
    .X(net321));
 sky130_fd_sc_hd__a21bo_1 c419 (.A1(net311),
    .A2(net215),
    .B1_N(net312),
    .X(net322));
 sky130_fd_sc_hd__a21bo_1 c420 (.A1(net810),
    .A2(net816),
    .B1_N(net224),
    .X(net323));
 sky130_fd_sc_hd__buf_1 c421 (.A(net690),
    .X(net324));
 sky130_fd_sc_hd__a21bo_1 c422 (.A1(net307),
    .A2(net301),
    .B1_N(net819),
    .X(net325));
 sky130_fd_sc_hd__xnor2_1 c423 (.A(net811),
    .B(net789),
    .Y(net326));
 sky130_fd_sc_hd__sdfbbn_2 c424 (.CLK_N(clknet_4_2_0_clk),
    .D(net844),
    .RESET_B(net799),
    .SCD(net322),
    .SCE(net209),
    .SET_B(net218),
    .Q(net328),
    .Q_N(net327));
 sky130_fd_sc_hd__a21bo_1 c425 (.A1(net799),
    .A2(net899),
    .B1_N(net327),
    .X(net329));
 sky130_fd_sc_hd__a21bo_1 c426 (.A1(net328),
    .A2(net792),
    .B1_N(net871),
    .X(net330));
 sky130_fd_sc_hd__dlymetal6s2s_1 c427 (.A(net777),
    .X(net331));
 sky130_fd_sc_hd__a41o_1 c428 (.A1(net329),
    .A2(net311),
    .A3(net898),
    .A4(net330),
    .B1(net906),
    .X(net332));
 sky130_fd_sc_hd__sdfbbn_2 c429 (.CLK_N(clknet_4_8_0_clk),
    .D(net844),
    .RESET_B(net898),
    .SCD(net205),
    .SCE(net332),
    .SET_B(net97),
    .Q(net334),
    .Q_N(net333));
 sky130_fd_sc_hd__clkbuf_1 c430 (.A(net690),
    .X(net335));
 sky130_fd_sc_hd__xnor2_2 c431 (.A(net331),
    .B(net334),
    .Y(net336));
 sky130_fd_sc_hd__a21bo_1 c432 (.A1(net222),
    .A2(net808),
    .B1_N(net928),
    .X(net337));
 sky130_fd_sc_hd__sdfsbp_2 c433 (.CLK(clknet_4_8_0_clk),
    .D(net196),
    .SCD(net218),
    .SCE(net336),
    .SET_B(net327),
    .Q(net339),
    .Q_N(net338));
 sky130_fd_sc_hd__a31o_1 c434 (.A1(net188),
    .A2(net335),
    .A3(net311),
    .B1(net924),
    .X(net340));
 sky130_fd_sc_hd__a21bo_2 c435 (.A1(net334),
    .A2(net305),
    .B1_N(net936),
    .X(net341));
 sky130_fd_sc_hd__a41o_1 c436 (.A1(net839),
    .A2(net318),
    .A3(net924),
    .A4(net901),
    .B1(net210),
    .X(net342));
 sky130_fd_sc_hd__mux4_2 c437 (.A0(net341),
    .A1(net312),
    .A2(net991),
    .A3(net910),
    .S0(net87),
    .S1(net923),
    .X(net343));
 sky130_fd_sc_hd__sdfbbp_1 c438 (.CLK(clknet_4_8_0_clk),
    .D(net335),
    .RESET_B(net327),
    .SCD(net341),
    .SCE(net923),
    .SET_B(net343),
    .Q(net345),
    .Q_N(net344));
 sky130_fd_sc_hd__a31o_1 c439 (.A1(net342),
    .A2(net341),
    .A3(net340),
    .B1(net923),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_2 c440 (.A(net646),
    .X(net868));
 sky130_fd_sc_hd__buf_1 c441 (.A(net645),
    .X(net347));
 sky130_fd_sc_hd__a21bo_1 c442 (.A1(net336),
    .A2(net868),
    .B1_N(net870),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_2 c443 (.A(net777),
    .X(net850));
 sky130_fd_sc_hd__a21bo_1 c444 (.A1(net326),
    .A2(net242),
    .B1_N(net344),
    .X(net349));
 sky130_fd_sc_hd__a21bo_1 c445 (.A1(net223),
    .A2(net348),
    .B1_N(clknet_1_0__leaf_net103),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_1 c446 (.A(net779),
    .X(net351));
 sky130_fd_sc_hd__sdfstp_1 c447 (.CLK(clknet_4_9_0_clk),
    .D(net236),
    .SCD(net321),
    .SCE(net227),
    .SET_B(net974),
    .Q(net352));
 sky130_fd_sc_hd__a21bo_1 c448 (.A1(clknet_1_1__leaf_net232),
    .A2(net798),
    .B1_N(net899),
    .X(net890));
 sky130_fd_sc_hd__mux4_2 c449 (.A0(net123),
    .A1(net798),
    .A2(net321),
    .A3(net96),
    .S0(net813),
    .S1(net348),
    .X(net353));
 sky130_fd_sc_hd__a41o_1 c450 (.A1(net352),
    .A2(net850),
    .A3(net301),
    .A4(net923),
    .B1(clknet_1_0__leaf_net350),
    .X(net354));
 sky130_fd_sc_hd__sdfbbn_1 c451 (.CLK_N(clknet_4_8_0_clk),
    .D(net332),
    .RESET_B(net981),
    .SCD(net336),
    .SCE(clknet_1_0__leaf_net354),
    .SET_B(net305),
    .Q(net356),
    .Q_N(net355));
 sky130_fd_sc_hd__a21bo_1 c452 (.A1(clknet_1_0__leaf_net230),
    .A2(net199),
    .B1_N(net349),
    .X(net357));
 sky130_fd_sc_hd__dlymetal6s2s_1 c453 (.A(net782),
    .X(net358));
 sky130_fd_sc_hd__a31o_1 c454 (.A1(net857),
    .A2(clknet_1_0__leaf_net354),
    .A3(net352),
    .B1(net692),
    .X(net359));
 sky130_fd_sc_hd__a21bo_1 c455 (.A1(clknet_1_0__leaf_net357),
    .A2(net347),
    .B1_N(net692),
    .X(net360));
 sky130_fd_sc_hd__sdfbbn_1 c456 (.CLK_N(clknet_4_9_0_clk),
    .D(net202),
    .RESET_B(clknet_1_0__leaf_net122),
    .SCD(net317),
    .SCE(net353),
    .SET_B(clknet_1_1__leaf_net354),
    .Q(net362),
    .Q_N(net361));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(clknet_1_1__leaf_net124),
    .A1(net352),
    .A2(clknet_1_0__leaf_net230),
    .A3(clknet_1_0__leaf_net354),
    .S0(clknet_1_1__leaf_net357),
    .S1(net687),
    .X(net363));
 sky130_fd_sc_hd__a41o_1 c458 (.A1(clknet_1_1__leaf_net360),
    .A2(clknet_1_0__leaf_net354),
    .A3(net352),
    .A4(net210),
    .B1(net236),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_2 c459 (.A(net968),
    .X(net365));
 sky130_fd_sc_hd__a41o_1 c460 (.A1(net73),
    .A2(net839),
    .A3(net365),
    .A4(clknet_1_0__leaf_net360),
    .B1(net714),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_1 c461 (.A(net779),
    .X(net367));
 sky130_fd_sc_hd__sdfbbp_1 c462 (.CLK(clknet_4_3_0_clk),
    .D(clknet_1_0__leaf_net366),
    .RESET_B(net309),
    .SCD(clknet_1_0__leaf_net233),
    .SCE(net262),
    .SET_B(clknet_1_0__leaf_net140),
    .Q(net369),
    .Q_N(net368));
 sky130_fd_sc_hd__mux4_1 c463 (.A0(net343),
    .A1(net817),
    .A2(net325),
    .A3(net318),
    .S0(net904),
    .S1(net228),
    .X(net370));
 sky130_fd_sc_hd__sdfbbn_1 c464 (.CLK_N(clknet_4_9_0_clk),
    .D(net325),
    .RESET_B(net853),
    .SCD(net227),
    .SCE(net312),
    .SET_B(net714),
    .Q(net372),
    .Q_N(net371));
 sky130_fd_sc_hd__a31o_1 c465 (.A1(clknet_1_1__leaf_net350),
    .A2(net820),
    .A3(clknet_1_0__leaf_net230),
    .B1(net20),
    .X(net373));
 sky130_fd_sc_hd__sdfstp_1 c466 (.CLK(clknet_4_3_0_clk),
    .D(net262),
    .SCD(net97),
    .SCE(net17),
    .SET_B(net917),
    .Q(net374));
 sky130_fd_sc_hd__mux4_1 c467 (.A0(net351),
    .A1(net365),
    .A2(net857),
    .A3(clknet_1_0__leaf_net124),
    .S0(clknet_1_0__leaf_net251),
    .S1(net248),
    .X(net375));
 sky130_fd_sc_hd__a41o_1 c468 (.A1(net8),
    .A2(net849),
    .A3(clknet_1_1__leaf_net268),
    .A4(net918),
    .B1(net722),
    .X(net376));
 sky130_fd_sc_hd__a41o_1 c469 (.A1(net198),
    .A2(net843),
    .A3(net799),
    .A4(net923),
    .B1(net714),
    .X(net377));
 sky130_fd_sc_hd__sdfstp_1 c470 (.CLK(clknet_4_3_0_clk),
    .D(net998),
    .SCD(net377),
    .SCE(net234),
    .SET_B(net318),
    .Q(net378));
 sky130_fd_sc_hd__sdfbbn_1 c471 (.CLK_N(clknet_4_3_0_clk),
    .D(net309),
    .RESET_B(net926),
    .SCD(net185),
    .SCE(clknet_1_1__leaf_net366),
    .SET_B(clknet_1_0__leaf_net376),
    .Q(net380),
    .Q_N(net379));
 sky130_fd_sc_hd__mux4_1 c472 (.A0(clknet_1_1__leaf_net124),
    .A1(net17),
    .A2(clknet_1_0__leaf_net270),
    .A3(net869),
    .S0(net20),
    .S1(net374),
    .X(net381));
 sky130_fd_sc_hd__a41o_1 c473 (.A1(clknet_1_0__leaf_net268),
    .A2(net829),
    .A3(net371),
    .A4(net20),
    .B1(net921),
    .X(net382));
 sky130_fd_sc_hd__a41o_1 c474 (.A1(net831),
    .A2(net918),
    .A3(clknet_1_0__leaf_net268),
    .A4(net714),
    .B1(net921),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 c475 (.A0(net926),
    .A1(net868),
    .A2(net214),
    .A3(clknet_1_0__leaf_net382),
    .S0(net998),
    .S1(net723),
    .X(net384));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(net384),
    .A1(net215),
    .A2(net374),
    .A3(clknet_1_0__leaf_net383),
    .S0(net870),
    .S1(clknet_1_1__leaf_net124),
    .X(net385));
 sky130_fd_sc_hd__a41o_1 c477 (.A1(clknet_1_1__leaf_net383),
    .A2(net147),
    .A3(net368),
    .A4(net792),
    .B1(net860),
    .X(net386));
 sky130_fd_sc_hd__a41o_1 c478 (.A1(net147),
    .A2(net228),
    .A3(net81),
    .A4(clknet_1_0__leaf_net386),
    .B1(clknet_1_0__leaf_net270),
    .X(net387));
 sky130_fd_sc_hd__a41o_1 c479 (.A1(net214),
    .A2(net81),
    .A3(clknet_1_0__leaf_net387),
    .A4(net898),
    .B1(net921),
    .X(net388));
 sky130_fd_sc_hd__sedfxbp_1 c480 (.CLK(clknet_4_3_0_clk),
    .D(clknet_1_0__leaf_net251),
    .DE(clknet_1_0__leaf_net695),
    .SCD(net722),
    .SCE(net921),
    .Q(net390),
    .Q_N(net389));
 sky130_fd_sc_hd__sdfbbp_1 c481 (.CLK(clknet_4_3_0_clk),
    .D(net983),
    .RESET_B(clknet_1_1__leaf_net387),
    .SCD(net389),
    .SCE(net952),
    .SET_B(net921),
    .Q(net392),
    .Q_N(net391));
 sky130_fd_sc_hd__a31o_1 c482 (.A1(net390),
    .A2(net868),
    .A3(net379),
    .B1(net921),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net248),
    .A1(clknet_1_1__leaf_net386),
    .A2(clknet_1_0__leaf_net382),
    .A3(net391),
    .S0(net916),
    .S1(net921),
    .X(net394));
 sky130_fd_sc_hd__mux4_2 c484 (.A0(net380),
    .A1(net38),
    .A2(net922),
    .A3(net157),
    .S0(net829),
    .S1(net713),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 c485 (.A0(net161),
    .A1(clknet_1_1__leaf_net134),
    .A2(net994),
    .A3(net952),
    .S0(net814),
    .S1(clknet_1_0__leaf_net863),
    .X(net396));
 sky130_fd_sc_hd__mux4_1 c486 (.A0(net158),
    .A1(net341),
    .A2(net795),
    .A3(clknet_1_1__leaf_net134),
    .S0(net159),
    .S1(clknet_1_1__leaf_net716),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 c487 (.A0(net193),
    .A1(net219),
    .A2(net157),
    .A3(net81),
    .S0(clknet_1_1__leaf_net290),
    .S1(net904),
    .X(net398));
 sky130_fd_sc_hd__mux4_1 c488 (.A0(net104),
    .A1(net158),
    .A2(net294),
    .A3(net688),
    .S0(clknet_1_0__leaf_net716),
    .S1(net726),
    .X(net399));
 sky130_fd_sc_hd__mux4_1 c489 (.A0(net81),
    .A1(net813),
    .A2(net69),
    .A3(net896),
    .S0(net277),
    .S1(clknet_1_1__leaf_net251),
    .X(net400));
 sky130_fd_sc_hd__mux4_1 c490 (.A0(net837),
    .A1(net396),
    .A2(net36),
    .A3(clknet_1_1__leaf_net251),
    .S0(net277),
    .S1(net713),
    .X(net401));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(net305),
    .A1(clknet_1_1__leaf_net129),
    .A2(net786),
    .A3(net166),
    .S0(net922),
    .S1(net713),
    .X(net402));
 sky130_fd_sc_hd__mux4_1 c492 (.A0(net312),
    .A1(net860),
    .A2(net872),
    .A3(net395),
    .S0(net837),
    .S1(net305),
    .X(net403));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(net185),
    .A1(net33),
    .A2(net318),
    .A3(clknet_1_0__leaf_net268),
    .S0(net845),
    .S1(net725),
    .X(net864));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(net813),
    .A1(net786),
    .A2(net277),
    .A3(net159),
    .S0(net151),
    .S1(net928),
    .X(net404));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(net848),
    .A1(net393),
    .A2(net276),
    .A3(net792),
    .S0(net726),
    .S1(net728),
    .X(net405));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(net378),
    .A1(clknet_1_1__leaf_net140),
    .A2(net829),
    .A3(net312),
    .S0(net697),
    .S1(net727),
    .X(net866));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net135),
    .A1(net157),
    .A2(net946),
    .A3(net795),
    .S0(net294),
    .S1(clknet_1_0__leaf_net290),
    .X(net406));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(net393),
    .A1(clknet_1_1__leaf_net251),
    .A2(net32),
    .A3(net846),
    .S0(clknet_1_1__leaf_net354),
    .S1(net318),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(net209),
    .A1(net37),
    .A2(net872),
    .A3(clknet_1_0__leaf_net866),
    .S0(net128),
    .S1(net345),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(net330),
    .A1(net403),
    .A2(net104),
    .A3(net971),
    .S0(net856),
    .S1(net810),
    .X(net409));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(net32),
    .A1(net408),
    .A2(net395),
    .A3(net725),
    .S0(net730),
    .S1(net731),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(net152),
    .A1(net406),
    .A2(net844),
    .A3(net185),
    .S0(net688),
    .S1(net731),
    .X(net411));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(net345),
    .A1(clknet_1_0__leaf_net866),
    .A2(net936),
    .A3(net166),
    .S0(net730),
    .S1(net731),
    .X(net412));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net318),
    .A1(net89),
    .A2(net994),
    .A3(net696),
    .S0(net730),
    .S1(net731),
    .X(net413));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(net405),
    .A1(net1001),
    .A2(clknet_1_1__leaf_net866),
    .A3(net786),
    .S0(net730),
    .S1(net732),
    .X(net414));
 sky130_fd_sc_hd__xnor2_4 c528 (.A(net843),
    .B(net817),
    .Y(net415));
 sky130_fd_sc_hd__xnor2_4 c529 (.A(net315),
    .B(net415),
    .Y(net416));
 sky130_fd_sc_hd__xnor2_1 c530 (.A(net73),
    .B(net797),
    .Y(net417));
 sky130_fd_sc_hd__buf_4 c531 (.A(net651),
    .X(net418));
 sky130_fd_sc_hd__xnor2_4 c532 (.A(net785),
    .B(net418),
    .Y(net419));
 sky130_fd_sc_hd__xnor2_4 c533 (.A(net792),
    .B(net842),
    .Y(net420));
 sky130_fd_sc_hd__xnor2_4 c534 (.A(net419),
    .B(net977),
    .Y(net894));
 sky130_fd_sc_hd__xnor2_4 c535 (.A(net302),
    .B(net200),
    .Y(net847));
 sky130_fd_sc_hd__buf_2 c536 (.A(net651),
    .X(net421));
 sky130_fd_sc_hd__a31o_2 c537 (.A1(net789),
    .A2(net194),
    .A3(net197),
    .B1(net418),
    .X(net422));
 sky130_fd_sc_hd__xnor2_2 c538 (.A(net817),
    .B(net421),
    .Y(net423));
 sky130_fd_sc_hd__xnor2_2 c539 (.A(net790),
    .B(net422),
    .Y(net424));
 sky130_fd_sc_hd__dlymetal6s2s_1 c540 (.A(net986),
    .X(net425));
 sky130_fd_sc_hd__xnor2_1 c541 (.A(net785),
    .B(net669),
    .Y(net426));
 sky130_fd_sc_hd__xnor2_2 c542 (.A(net303),
    .B(net306),
    .Y(net427));
 sky130_fd_sc_hd__xnor2_4 c543 (.A(net828),
    .B(net416),
    .Y(net428));
 sky130_fd_sc_hd__a31o_1 c544 (.A1(net427),
    .A2(net421),
    .A3(net319),
    .B1(net300),
    .X(net429));
 sky130_fd_sc_hd__a31o_1 c545 (.A1(net418),
    .A2(net429),
    .A3(net420),
    .B1(net314),
    .X(net430));
 sky130_fd_sc_hd__xnor2_1 c546 (.A(net420),
    .B(net644),
    .Y(net431));
 sky130_fd_sc_hd__xnor2_1 c547 (.A(net428),
    .B(net678),
    .Y(net432));
 sky130_fd_sc_hd__xnor2_1 c548 (.A(net426),
    .B(net421),
    .Y(net433));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(net432),
    .A1(net424),
    .A2(net431),
    .A3(net425),
    .S0(net419),
    .S1(net421),
    .X(net434));
 sky130_fd_sc_hd__xnor2_1 c550 (.A(net816),
    .B(net428),
    .Y(net435));
 sky130_fd_sc_hd__a21bo_1 c551 (.A1(net435),
    .A2(net224),
    .B1_N(net910),
    .X(net436));
 sky130_fd_sc_hd__mux4_1 c552 (.A0(net331),
    .A1(net899),
    .A2(net213),
    .A3(net900),
    .S0(net923),
    .S1(clknet_1_0__leaf_net733),
    .X(net437));
 sky130_fd_sc_hd__a21bo_1 c553 (.A1(net426),
    .A2(net337),
    .B1_N(clknet_1_1__leaf_net733),
    .X(net438));
 sky130_fd_sc_hd__xnor2_1 c554 (.A(net87),
    .B(clknet_1_0__leaf_net437),
    .Y(net439));
 sky130_fd_sc_hd__a21bo_1 c555 (.A1(net842),
    .A2(net894),
    .B1_N(clknet_1_1__leaf_net439),
    .X(net440));
 sky130_fd_sc_hd__buf_1 c556 (.A(net706),
    .X(net441));
 sky130_fd_sc_hd__a21bo_1 c557 (.A1(net421),
    .A2(net441),
    .B1_N(net819),
    .X(net442));
 sky130_fd_sc_hd__a21bo_1 c558 (.A1(net320),
    .A2(clknet_1_0__leaf_net437),
    .B1_N(net324),
    .X(net443));
 sky130_fd_sc_hd__xnor2_1 c559 (.A(net794),
    .B(net415),
    .Y(net444));
 sky130_fd_sc_hd__a31o_1 c560 (.A1(net442),
    .A2(net324),
    .A3(net191),
    .B1(net928),
    .X(net445));
 sky130_fd_sc_hd__a21bo_2 c561 (.A1(net218),
    .A2(net910),
    .B1_N(net785),
    .X(net446));
 sky130_fd_sc_hd__mux4_1 c562 (.A0(net803),
    .A1(net418),
    .A2(net446),
    .A3(net419),
    .S0(net89),
    .S1(net415),
    .X(net447));
 sky130_fd_sc_hd__a21bo_1 c563 (.A1(net445),
    .A2(net442),
    .B1_N(clknet_1_0__leaf_net733),
    .X(net448));
 sky130_fd_sc_hd__xnor2_4 c564 (.A(net416),
    .B(net692),
    .Y(net449));
 sky130_fd_sc_hd__xnor2_1 c565 (.A(clknet_1_1__leaf_net437),
    .B(net445),
    .Y(net450));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(net450),
    .A1(net222),
    .A2(net333),
    .A3(net446),
    .S0(net449),
    .S1(clknet_1_0__leaf_net448),
    .X(net451));
 sky130_fd_sc_hd__a21bo_2 c567 (.A1(net444),
    .A2(net919),
    .B1_N(net923),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_1 c568 (.A(net706),
    .X(net452));
 sky130_fd_sc_hd__xnor2_2 c569 (.A(net324),
    .B(net213),
    .Y(net453));
 sky130_fd_sc_hd__a21bo_1 c570 (.A1(net452),
    .A2(net445),
    .B1_N(net447),
    .X(net454));
 sky130_fd_sc_hd__xnor2_1 c571 (.A(net337),
    .B(clknet_1_1__leaf_net437),
    .Y(net455));
 sky130_fd_sc_hd__a31o_1 c572 (.A1(net447),
    .A2(clknet_1_1__leaf_net122),
    .A3(net321),
    .B1(net427),
    .X(net456));
 sky130_fd_sc_hd__a21bo_1 c573 (.A1(net242),
    .A2(net818),
    .B1_N(clknet_1_0__leaf_net239),
    .X(net457));
 sky130_fd_sc_hd__a21bo_1 c574 (.A1(net453),
    .A2(net928),
    .B1_N(net207),
    .X(net458));
 sky130_fd_sc_hd__a31o_1 c575 (.A1(net417),
    .A2(net841),
    .A3(net429),
    .B1(net818),
    .X(net459));
 sky130_fd_sc_hd__sedfxbp_2 c576 (.CLK(clknet_4_9_0_clk),
    .D(net348),
    .DE(net73),
    .SCD(net853),
    .SCE(net669),
    .Q(net461),
    .Q_N(net460));
 sky130_fd_sc_hd__sedfxtp_1 c577 (.CLK(clknet_4_9_0_clk),
    .D(net96),
    .DE(net234),
    .SCD(clknet_1_0__leaf_net443),
    .SCE(net454),
    .Q(net462));
 sky130_fd_sc_hd__a31o_1 c578 (.A1(net429),
    .A2(clknet_1_0__leaf_net457),
    .A3(net840),
    .B1(clknet_1_1__leaf_net120),
    .X(net463));
 sky130_fd_sc_hd__a31o_1 c579 (.A1(net415),
    .A2(net334),
    .A3(net73),
    .B1(net210),
    .X(net464));
 sky130_fd_sc_hd__a31o_1 c580 (.A1(net825),
    .A2(clknet_1_0__leaf_net116),
    .A3(net415),
    .B1(net453),
    .X(net465));
 sky130_fd_sc_hd__a41o_1 c581 (.A1(net367),
    .A2(net321),
    .A3(net847),
    .A4(net850),
    .B1(clknet_1_1__leaf_net465),
    .X(net466));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(net459),
    .A1(net456),
    .A2(clknet_1_0__leaf_net890),
    .A3(clknet_1_1__leaf_net465),
    .S0(net789),
    .S1(net785),
    .X(net467));
 sky130_fd_sc_hd__mux4_1 c583 (.A0(net231),
    .A1(clknet_1_0__leaf_net116),
    .A2(net462),
    .A3(net73),
    .S0(net901),
    .S1(net418),
    .X(net468));
 sky130_fd_sc_hd__a31o_1 c584 (.A1(clknet_1_1__leaf_net117),
    .A2(net453),
    .A3(clknet_1_0__leaf_net465),
    .B1(net923),
    .X(net469));
 sky130_fd_sc_hd__a41o_1 c585 (.A1(clknet_1_1__leaf_net116),
    .A2(net328),
    .A3(net855),
    .A4(net417),
    .B1(clknet_1_0__leaf_net734),
    .X(net470));
 sky130_fd_sc_hd__a31o_1 c586 (.A1(net470),
    .A2(clknet_1_0__leaf_net465),
    .A3(net89),
    .B1(net210),
    .X(net471));
 sky130_fd_sc_hd__a21bo_1 c587 (.A1(net210),
    .A2(clknet_1_0__leaf_net471),
    .B1_N(clknet_1_0__leaf_net463),
    .X(net472));
 sky130_fd_sc_hd__a31o_1 c588 (.A1(net441),
    .A2(clknet_1_0__leaf_net472),
    .A3(net203),
    .B1(clknet_1_0__leaf_net465),
    .X(net473));
 sky130_fd_sc_hd__sdfbbn_1 c589 (.CLK_N(clknet_4_9_0_clk),
    .D(net454),
    .RESET_B(net347),
    .SCD(clknet_1_1__leaf_net472),
    .SCE(net361),
    .SET_B(clknet_1_0__leaf_net465),
    .Q(net475),
    .Q_N(net474));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(net451),
    .A1(net459),
    .A2(net415),
    .A3(net474),
    .S0(net898),
    .S1(clknet_1_1__leaf_net465),
    .X(net476));
 sky130_fd_sc_hd__a41o_1 c591 (.A1(net213),
    .A2(net356),
    .A3(clknet_1_1__leaf_net457),
    .A4(clknet_1_1__leaf_net465),
    .B1(clknet_1_0__leaf_net694),
    .X(net477));
 sky130_fd_sc_hd__a41o_1 c592 (.A1(net458),
    .A2(net365),
    .A3(clknet_1_0__leaf_net469),
    .A4(clknet_1_0__leaf_net455),
    .B1(clknet_1_0__leaf_net465),
    .X(net478));
 sky130_fd_sc_hd__a41o_1 c593 (.A1(clknet_1_1__leaf_net469),
    .A2(clknet_1_0__leaf_net478),
    .A3(net454),
    .A4(net358),
    .B1(clknet_1_1__leaf_net734),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c594 (.A0(net802),
    .A1(clknet_1_1__leaf_net142),
    .A2(net924),
    .A3(net301),
    .S0(clknet_1_1__leaf_net268),
    .S1(net683),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c595 (.A0(clknet_1_0__leaf_net448),
    .A1(net787),
    .A2(net200),
    .A3(net424),
    .S0(net906),
    .S1(net713),
    .X(net481));
 sky130_fd_sc_hd__a41o_1 c596 (.A1(net17),
    .A2(net908),
    .A3(net924),
    .A4(clknet_1_1__leaf_net270),
    .B1(net1009),
    .X(net482));
 sky130_fd_sc_hd__mux4_1 c597 (.A0(net207),
    .A1(net480),
    .A2(clknet_1_1__leaf_net103),
    .A3(net365),
    .S0(net723),
    .S1(net725),
    .X(net483));
 sky130_fd_sc_hd__a41o_1 c598 (.A1(net227),
    .A2(net89),
    .A3(net810),
    .A4(net419),
    .B1(net831),
    .X(net484));
 sky130_fd_sc_hd__mux4_2 c599 (.A0(clknet_1_1__leaf_net382),
    .A1(net417),
    .A2(clknet_1_1__leaf_net448),
    .A3(net328),
    .S0(net321),
    .S1(net17),
    .X(net485));
 sky130_fd_sc_hd__sdfbbn_1 c600 (.CLK_N(clknet_4_14_0_clk),
    .D(net464),
    .RESET_B(clknet_1_1__leaf_net233),
    .SCD(net793),
    .SCE(net929),
    .SET_B(clknet_1_0__leaf_net485),
    .Q(net487),
    .Q_N(net486));
 sky130_fd_sc_hd__mux4_1 c601 (.A0(net213),
    .A1(net328),
    .A2(net484),
    .A3(net894),
    .S0(net898),
    .S1(clknet_1_1__leaf_net268),
    .X(net488));
 sky130_fd_sc_hd__a41o_1 c602 (.A1(net362),
    .A2(net819),
    .A3(net944),
    .A4(clknet_1_1__leaf_net268),
    .B1(net904),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(clknet_1_1__leaf_net270),
    .A1(clknet_1_0__leaf_net489),
    .A2(net464),
    .A3(net808),
    .S0(clknet_1_0__leaf_net465),
    .S1(net724),
    .X(net893));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(net301),
    .A1(net813),
    .A2(net211),
    .A3(net227),
    .S0(net855),
    .S1(clknet_1_1__leaf_net489),
    .X(net490));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(clknet_1_1__leaf_net112),
    .A1(net794),
    .A2(net227),
    .A3(net916),
    .S0(clknet_1_1__leaf_net268),
    .S1(net725),
    .X(net491));
 sky130_fd_sc_hd__a41o_1 c606 (.A1(net831),
    .A2(clknet_1_0__leaf_net890),
    .A3(net328),
    .B1(clknet_1_0__leaf_net735),
    .X(net492));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(net483),
    .A1(net201),
    .A2(net362),
    .A3(net484),
    .S0(net788),
    .S1(clknet_1_0__leaf_net122),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net431),
    .A1(net904),
    .A2(net789),
    .A3(net923),
    .S0(net672),
    .S1(net724),
    .X(net494));
 sky130_fd_sc_hd__a41o_1 c609 (.A1(net419),
    .A2(net475),
    .A3(net848),
    .A4(clknet_1_1__leaf_net112),
    .B1(clknet_1_1__leaf_net268),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c610 (.A0(net808),
    .A1(clknet_1_1__leaf_net140),
    .A2(net916),
    .A3(net911),
    .S0(net937),
    .S1(net921),
    .X(net862));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net372),
    .A1(net495),
    .A2(net102),
    .A3(clknet_1_1__leaf_net376),
    .S0(clknet_1_1__leaf_net270),
    .S1(net852),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(net321),
    .A1(net853),
    .A2(net428),
    .A3(net924),
    .S0(net918),
    .S1(net994),
    .X(net497));
 sky130_fd_sc_hd__a41o_1 c613 (.A1(net418),
    .A2(net236),
    .A3(net8),
    .A4(net929),
    .B1(net965),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(net798),
    .A1(net219),
    .A2(net810),
    .A3(net17),
    .S0(net794),
    .S1(net737),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net8),
    .A1(net207),
    .A2(net17),
    .A3(clknet_1_0__leaf_net489),
    .S0(net700),
    .S1(net738),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c616 (.A0(net812),
    .A1(clknet_1_0__leaf_net468),
    .A2(net826),
    .A3(net295),
    .S0(net946),
    .S1(net128),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(net104),
    .A1(net908),
    .A2(net108),
    .A3(net906),
    .S0(net785),
    .S1(net669),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(net848),
    .A1(net284),
    .A2(net845),
    .A3(net141),
    .S0(net62),
    .S1(net718),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c619 (.A0(net428),
    .A1(net462),
    .A2(net936),
    .A3(net283),
    .S0(clknet_1_1__leaf_net120),
    .S1(clknet_1_1__leaf_net140),
    .X(net504));
 sky130_fd_sc_hd__mux4_2 c62 (.A0(net824),
    .A1(net833),
    .A2(net796),
    .A3(net823),
    .S0(net812),
    .S1(net834),
    .X(net0));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net402),
    .A1(net104),
    .A2(net930),
    .A3(net219),
    .S0(net986),
    .S1(net725),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(net141),
    .A1(net994),
    .A2(net414),
    .A3(net786),
    .S0(net333),
    .S1(net731),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(net424),
    .A1(net300),
    .A2(net916),
    .A3(net159),
    .S0(net644),
    .S1(net854),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(net146),
    .A1(net159),
    .A2(net413),
    .A3(net69),
    .S0(net848),
    .S1(net952),
    .X(net508));
 sky130_fd_sc_hd__mux4_1 c624 (.A0(net102),
    .A1(net288),
    .A2(net369),
    .A3(clknet_1_1__leaf_net268),
    .S0(net1009),
    .S1(net275),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net980),
    .A1(net504),
    .A2(clknet_1_0__leaf_net376),
    .A3(net300),
    .S0(net1007),
    .S1(net725),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net843),
    .A1(clknet_1_1__leaf_net290),
    .A2(net812),
    .A3(net288),
    .S0(clknet_1_0__leaf_net412),
    .S1(clknet_1_1__leaf_net478),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(net219),
    .A1(net369),
    .A2(clknet_1_0__leaf_net412),
    .A3(net851),
    .S0(net994),
    .S1(net729),
    .X(net512));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net503),
    .A1(net644),
    .A2(clknet_1_1__leaf_net140),
    .A3(net845),
    .S0(net847),
    .S1(clknet_1_0__leaf_net268),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(net277),
    .A1(net108),
    .A2(net812),
    .A3(clknet_1_1__leaf_net103),
    .S0(net428),
    .S1(net945),
    .X(net514));
 sky130_fd_sc_hd__mux4_2 c63 (.A0(net833),
    .A1(net827),
    .A2(net835),
    .A3(net830),
    .S0(net840),
    .S1(net829),
    .X(net852));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net449),
    .A1(clknet_1_1__leaf_net463),
    .A2(net904),
    .A3(net786),
    .S0(net906),
    .S1(net739),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net494),
    .A1(net484),
    .A2(net852),
    .A3(net894),
    .S0(net813),
    .S1(net726),
    .X(net516));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net89),
    .A1(net166),
    .A2(net904),
    .A3(net812),
    .S0(net276),
    .S1(clknet_1_0__leaf_net515),
    .X(net517));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(net488),
    .A1(net449),
    .A2(clknet_1_1__leaf_net142),
    .A3(clknet_1_1__leaf_net120),
    .S0(net873),
    .S1(net742),
    .X(net518));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net276),
    .A1(net484),
    .A2(net996),
    .A3(net449),
    .S0(clknet_1_0__leaf_net282),
    .S1(net741),
    .X(net519));
 sky130_fd_sc_hd__mux4_2 c635 (.A0(net514),
    .A1(net916),
    .A2(net792),
    .A3(net333),
    .S0(net918),
    .S1(net705),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net516),
    .A1(net785),
    .A2(clknet_1_1__leaf_net468),
    .A3(clknet_1_0__leaf_net493),
    .S0(clknet_1_1__leaf_net735),
    .S1(net743),
    .X(net521));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net145),
    .A1(net1001),
    .A2(clknet_1_0__leaf_net493),
    .A3(net680),
    .S0(net723),
    .S1(net744),
    .X(net522));
 sky130_fd_sc_hd__mux4_2 c64 (.A0(net819),
    .A1(net829),
    .A2(net840),
    .A3(net839),
    .S0(net825),
    .S1(net0),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c65 (.A0(net822),
    .A1(net804),
    .A2(net1013),
    .A3(net795),
    .S0(net824),
    .S1(net819),
    .X(net2));
 sky130_fd_sc_hd__xnor2_4 c66 (.A(net829),
    .B(net832),
    .Y(net3));
 sky130_fd_sc_hd__a21bo_1 c660 (.A1(net313),
    .A2(net433),
    .B1_N(net900),
    .X(net523));
 sky130_fd_sc_hd__xnor2_1 c661 (.A(net828),
    .B(net898),
    .Y(net524));
 sky130_fd_sc_hd__xnor2_2 c662 (.A(net828),
    .B(net523),
    .Y(net525));
 sky130_fd_sc_hd__xnor2_1 c663 (.A(net194),
    .B(net900),
    .Y(net526));
 sky130_fd_sc_hd__xnor2_2 c664 (.A(net310),
    .B(net919),
    .Y(net527));
 sky130_fd_sc_hd__xnor2_2 c665 (.A(net420),
    .B(net942),
    .Y(net528));
 sky130_fd_sc_hd__xnor2_1 c666 (.A(net433),
    .B(net425),
    .Y(net529));
 sky130_fd_sc_hd__a21bo_1 c667 (.A1(net527),
    .A2(net306),
    .B1_N(net912),
    .X(net530));
 sky130_fd_sc_hd__xnor2_1 c668 (.A(net523),
    .B(net197),
    .Y(net531));
 sky130_fd_sc_hd__buf_1 c669 (.A(net686),
    .X(net532));
 sky130_fd_sc_hd__xnor2_4 c67 (.A(net823),
    .B(net822),
    .Y(net4));
 sky130_fd_sc_hd__buf_1 c670 (.A(net699),
    .X(net533));
 sky130_fd_sc_hd__xnor2_1 c671 (.A(net197),
    .B(net930),
    .Y(net534));
 sky130_fd_sc_hd__a21bo_1 c672 (.A1(net531),
    .A2(net525),
    .B1_N(net529),
    .X(net535));
 sky130_fd_sc_hd__mux4_1 c673 (.A0(net530),
    .A1(net899),
    .A2(net527),
    .A3(net528),
    .S0(net197),
    .S1(net919),
    .X(net536));
 sky130_fd_sc_hd__xnor2_1 c674 (.A(net529),
    .B(net532),
    .Y(net537));
 sky130_fd_sc_hd__dlymetal6s2s_1 c675 (.A(net698),
    .X(net538));
 sky130_fd_sc_hd__a21bo_1 c676 (.A1(net797),
    .A2(net943),
    .B1_N(net537),
    .X(net539));
 sky130_fd_sc_hd__buf_1 c677 (.A(net685),
    .X(net540));
 sky130_fd_sc_hd__a21bo_1 c678 (.A1(net536),
    .A2(net527),
    .B1_N(net538),
    .X(net541));
 sky130_fd_sc_hd__buf_2 c679 (.A(net698),
    .X(net542));
 sky130_fd_sc_hd__xnor2_4 c68 (.A(net1013),
    .B(net4),
    .Y(net5));
 sky130_fd_sc_hd__a21bo_1 c680 (.A1(net537),
    .A2(net194),
    .B1_N(net542),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_2 c681 (.A(net686),
    .X(net544));
 sky130_fd_sc_hd__a31o_1 c682 (.A1(net528),
    .A2(clknet_1_0__leaf_net439),
    .A3(net533),
    .B1(net340),
    .X(net545));
 sky130_fd_sc_hd__a41o_1 c683 (.A1(clknet_1_1__leaf_net545),
    .A2(net425),
    .A3(net899),
    .A4(clknet_1_0__leaf_net103),
    .B1(net790),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_1 c684 (.A(net685),
    .X(net547));
 sky130_fd_sc_hd__a31o_1 c685 (.A1(net900),
    .A2(net423),
    .A3(net899),
    .B1(clknet_1_0__leaf_net438),
    .X(net548));
 sky130_fd_sc_hd__a31o_1 c686 (.A1(net346),
    .A2(net422),
    .A3(net924),
    .B1(net446),
    .X(net549));
 sky130_fd_sc_hd__a31o_1 c687 (.A1(net533),
    .A2(net539),
    .A3(net446),
    .B1(clknet_1_0__leaf_net103),
    .X(net550));
 sky130_fd_sc_hd__a31o_1 c688 (.A1(clknet_1_1__leaf_net550),
    .A2(net544),
    .A3(net446),
    .B1(net924),
    .X(net551));
 sky130_fd_sc_hd__sdfbbp_1 c689 (.CLK(clknet_4_10_0_clk),
    .D(net436),
    .RESET_B(net346),
    .SCD(net542),
    .SCE(net544),
    .SET_B(net1013),
    .Q(net553),
    .Q_N(net552));
 sky130_fd_sc_hd__a21bo_4 c69 (.A1(net805),
    .A2(net844),
    .B1_N(net833),
    .X(net6));
 sky130_fd_sc_hd__a31o_1 c690 (.A1(net540),
    .A2(net924),
    .A3(net927),
    .B1(net984),
    .X(net554));
 sky130_fd_sc_hd__a31o_1 c691 (.A1(net217),
    .A2(net542),
    .A3(net801),
    .B1(net552),
    .X(net555));
 sky130_fd_sc_hd__a21bo_1 c692 (.A1(net217),
    .A2(net552),
    .B1_N(net692),
    .X(net556));
 sky130_fd_sc_hd__a31o_2 c693 (.A1(net422),
    .A2(net539),
    .A3(net553),
    .B1(net818),
    .X(net557));
 sky130_fd_sc_hd__mux4_1 c694 (.A0(net340),
    .A1(net331),
    .A2(net557),
    .A3(net538),
    .S0(net818),
    .S1(net927),
    .X(net558));
 sky130_fd_sc_hd__a31o_1 c695 (.A1(clknet_1_0__leaf_net440),
    .A2(net534),
    .A3(net553),
    .B1(net538),
    .X(net559));
 sky130_fd_sc_hd__a31o_1 c696 (.A1(net425),
    .A2(net797),
    .A3(net317),
    .B1(clknet_1_0__leaf_net550),
    .X(net560));
 sky130_fd_sc_hd__sdfbbn_1 c697 (.CLK_N(clknet_4_10_0_clk),
    .D(net797),
    .RESET_B(net422),
    .SCD(net530),
    .SCE(net900),
    .SET_B(net557),
    .Q(net562),
    .Q_N(net561));
 sky130_fd_sc_hd__a31o_1 c698 (.A1(net534),
    .A2(net919),
    .A3(net533),
    .B1(net982),
    .X(net563));
 sky130_fd_sc_hd__sdfbbn_1 c699 (.CLK_N(clknet_4_10_0_clk),
    .D(net790),
    .RESET_B(net895),
    .SCD(clknet_1_0__leaf_net548),
    .SCE(clknet_1_0__leaf_net455),
    .SET_B(net528),
    .Q(net565),
    .Q_N(net564));
 sky130_fd_sc_hd__xnor2_4 c70 (.A(net821),
    .B(net824),
    .Y(net7));
 sky130_fd_sc_hd__sdfbbp_1 c700 (.CLK(clknet_4_10_0_clk),
    .D(net895),
    .RESET_B(net554),
    .SCD(net564),
    .SCE(net967),
    .SET_B(net982),
    .Q(net567),
    .Q_N(net566));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(net801),
    .A1(clknet_1_1__leaf_net440),
    .A2(net900),
    .A3(net566),
    .S0(net895),
    .S1(net984),
    .X(net568));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net224),
    .A1(net543),
    .A2(net539),
    .A3(net895),
    .S0(net211),
    .S1(net749),
    .X(net569));
 sky130_fd_sc_hd__sdfbbn_1 c703 (.CLK_N(clknet_4_10_0_clk),
    .D(net555),
    .RESET_B(net436),
    .SCD(net895),
    .SCE(net561),
    .SET_B(clknet_1_0__leaf_net750),
    .Q(net571),
    .Q_N(net570));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net356),
    .A1(net906),
    .A2(clknet_1_1__leaf_net465),
    .A3(net942),
    .S0(net787),
    .S1(net842),
    .X(net572));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(net801),
    .A1(clknet_1_1__leaf_net114),
    .A2(clknet_1_1__leaf_net465),
    .A3(clknet_1_0__leaf_net103),
    .S0(net432),
    .S1(net901),
    .X(net573));
 sky130_fd_sc_hd__sdfbbn_1 c706 (.CLK_N(clknet_4_10_0_clk),
    .D(net978),
    .RESET_B(net906),
    .SCD(net205),
    .SCE(net841),
    .SET_B(clknet_1_0__leaf_net551),
    .Q(net575),
    .Q_N(net574));
 sky130_fd_sc_hd__mux4_1 c707 (.A0(net205),
    .A1(net962),
    .A2(clknet_1_1__leaf_net239),
    .A3(net575),
    .S0(net787),
    .S1(clknet_1_1__leaf_net560),
    .X(net576));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(net538),
    .A1(clknet_1_1__leaf_net443),
    .A2(net542),
    .A3(net205),
    .S0(clknet_1_1__leaf_net438),
    .S1(clknet_1_0__leaf_net455),
    .X(net577));
 sky130_fd_sc_hd__sdfbbp_1 c709 (.CLK(clknet_4_11_0_clk),
    .D(net840),
    .RESET_B(net1010),
    .SCD(net538),
    .SCE(net535),
    .SET_B(net964),
    .Q(net579),
    .Q_N(net578));
 sky130_fd_sc_hd__xnor2_4 c71 (.A(net839),
    .B(net815),
    .Y(net8));
 sky130_fd_sc_hd__sdfbbn_1 c710 (.CLK_N(clknet_4_11_0_clk),
    .D(clknet_1_1__leaf_net239),
    .RESET_B(net838),
    .SCD(net317),
    .SCE(clknet_1_1__leaf_net122),
    .SET_B(net895),
    .Q(net581),
    .Q_N(net580));
 sky130_fd_sc_hd__a41o_1 c711 (.A1(net432),
    .A2(net477),
    .A3(clknet_1_0__leaf_net239),
    .A4(net317),
    .B1(net423),
    .X(net582));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net530),
    .A1(net547),
    .A2(net793),
    .A3(clknet_1_1__leaf_net694),
    .S0(clknet_1_0__leaf_net750),
    .S1(clknet_1_0__leaf_net751),
    .X(net583));
 sky130_fd_sc_hd__sdfbbn_1 c713 (.CLK_N(clknet_4_10_0_clk),
    .D(net446),
    .RESET_B(net802),
    .SCD(net841),
    .SCE(net557),
    .SET_B(net749),
    .Q(net585),
    .Q_N(net584));
 sky130_fd_sc_hd__sdfbbp_1 c714 (.CLK(clknet_4_14_0_clk),
    .D(net317),
    .RESET_B(net962),
    .SCD(net563),
    .SCE(net930),
    .SET_B(clknet_1_1__leaf_net752),
    .Q(net587),
    .Q_N(net586));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(clknet_1_0__leaf_net572),
    .A1(net535),
    .A2(net355),
    .A3(net930),
    .S0(clknet_1_0__leaf_net103),
    .S1(net552),
    .X(net588));
 sky130_fd_sc_hd__sdfbbn_1 c716 (.CLK_N(clknet_4_11_0_clk),
    .D(clknet_1_0__leaf_net438),
    .RESET_B(net525),
    .SCD(net895),
    .SCE(clknet_1_1__leaf_net572),
    .SET_B(net787),
    .Q(net590),
    .Q_N(net589));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net583),
    .A1(net927),
    .A2(net580),
    .A3(net928),
    .S0(net895),
    .S1(net201),
    .X(net591));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(net793),
    .A1(net585),
    .A2(clknet_1_1__leaf_net239),
    .A3(net901),
    .S0(net924),
    .S1(net460),
    .X(net592));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net553),
    .A1(net584),
    .A2(clknet_1_0__leaf_net354),
    .A3(net895),
    .S0(clknet_1_0__leaf_net750),
    .S1(net756),
    .X(net593));
 sky130_fd_sc_hd__xnor2_4 c72 (.A(net5),
    .B(net3),
    .Y(net9));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(clknet_1_0__leaf_net582),
    .A1(net581),
    .A2(clknet_1_1__leaf_net592),
    .A3(net906),
    .S0(clknet_1_0__leaf_net103),
    .S1(net755),
    .X(net594));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net899),
    .A1(net589),
    .A2(net201),
    .A3(net543),
    .S0(net820),
    .S1(net666),
    .X(net595));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net820),
    .A1(net578),
    .A2(net544),
    .A3(net919),
    .S0(net789),
    .S1(clknet_1_1__leaf_net751),
    .X(net596));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net838),
    .A1(net567),
    .A2(net840),
    .A3(clknet_1_1__leaf_net122),
    .S0(net446),
    .S1(net757),
    .X(net597));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(clknet_1_1__leaf_net551),
    .A1(clknet_1_0__leaf_net592),
    .A2(net525),
    .A3(net841),
    .S0(clknet_1_1__leaf_net597),
    .S1(net754),
    .X(net598));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net841),
    .A1(clknet_1_1__leaf_net582),
    .A2(clknet_1_0__leaf_net465),
    .A3(net317),
    .S0(net574),
    .S1(net758),
    .X(net599));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net547),
    .A1(clknet_1_1__leaf_net122),
    .A2(net427),
    .A3(clknet_1_1__leaf_net268),
    .S0(net708),
    .S1(net759),
    .X(net600));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net562),
    .A1(net571),
    .A2(clknet_1_1__leaf_net455),
    .A3(net228),
    .S0(clknet_1_0__leaf_net596),
    .S1(net784),
    .X(net601));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(clknet_1_1__leaf_net103),
    .A1(clknet_1_1__leaf_net455),
    .A2(net787),
    .A3(clknet_1_1__leaf_net485),
    .S0(net700),
    .S1(net759),
    .X(net602));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(net944),
    .A1(net200),
    .A2(net946),
    .A3(net842),
    .S0(net963),
    .S1(clknet_1_0__leaf_net478),
    .X(net603));
 sky130_fd_sc_hd__xnor2_4 c73 (.A(net806),
    .B(net821),
    .Y(net10));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(clknet_1_1__leaf_net136),
    .A1(net203),
    .A2(net586),
    .A3(net228),
    .S0(clknet_1_1__leaf_net103),
    .S1(net898),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net929),
    .A1(net544),
    .A2(clknet_1_1__leaf_net596),
    .A3(net557),
    .S0(net1006),
    .S1(net358),
    .X(net605));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(net423),
    .A1(net542),
    .A2(net788),
    .A3(net929),
    .S0(clknet_1_1__leaf_net750),
    .S1(net753),
    .X(net606));
 sky130_fd_sc_hd__mux4_2 c733 (.A0(net842),
    .A1(net793),
    .A2(net789),
    .A3(net487),
    .S0(net927),
    .S1(net703),
    .X(net607));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(net587),
    .A1(net487),
    .A2(net203),
    .A3(net820),
    .S0(net228),
    .S1(net787),
    .X(net608));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(clknet_1_1__leaf_net127),
    .A1(net570),
    .A2(net544),
    .A3(net8),
    .S0(net929),
    .S1(clknet_1_0__leaf_net752),
    .X(net609));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(net8),
    .A1(net787),
    .A2(net543),
    .A3(net901),
    .S0(net753),
    .S1(net761),
    .X(net610));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net557),
    .A1(clknet_1_1__leaf_net471),
    .A2(net579),
    .A3(net901),
    .S0(net8),
    .S1(net921),
    .X(net611));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net901),
    .A1(net802),
    .A2(net788),
    .A3(net607),
    .S0(net720),
    .S1(net761),
    .X(net612));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(net985),
    .A1(net600),
    .A2(net544),
    .A3(net8),
    .S0(net665),
    .S1(net713),
    .X(net613));
 sky130_fd_sc_hd__a21bo_4 c74 (.A1(net10),
    .A2(net820),
    .B1_N(net837),
    .X(net11));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(net963),
    .A1(net563),
    .A2(net543),
    .A3(net918),
    .S0(net677),
    .S1(net993),
    .X(net614));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(clknet_1_0__leaf_net597),
    .A1(net373),
    .A2(clknet_1_0__leaf_net485),
    .A3(net936),
    .S0(net929),
    .S1(net8),
    .X(net615));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(net211),
    .A1(net1006),
    .A2(net85),
    .A3(net542),
    .S0(net895),
    .S1(net973),
    .X(net616));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(net606),
    .A1(net842),
    .A2(net607),
    .A3(clknet_1_1__leaf_net750),
    .S0(net754),
    .S1(net761),
    .X(net617));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(net500),
    .A1(net595),
    .A2(clknet_1_0__leaf_net617),
    .A3(net802),
    .S0(net929),
    .S1(net708),
    .X(net618));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(clknet_1_0__leaf_net465),
    .A1(net543),
    .A2(net590),
    .A3(net924),
    .S0(net19),
    .S1(net761),
    .X(net619));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net228),
    .A1(net618),
    .A2(clknet_1_0__leaf_net619),
    .A3(net333),
    .S0(net195),
    .S1(net486),
    .X(net620));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(net927),
    .A1(net358),
    .A2(net612),
    .A3(net228),
    .S0(clknet_1_1__leaf_net619),
    .S1(net836),
    .X(net621));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net365),
    .A1(net989),
    .A2(net275),
    .A3(net1007),
    .S0(net745),
    .S1(net993),
    .X(net622));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net610),
    .A1(net961),
    .A2(clknet_1_1__leaf_net282),
    .A3(clknet_1_1__leaf_net412),
    .S0(clknet_1_1__leaf_net103),
    .S1(net768),
    .X(net623));
 sky130_fd_sc_hd__xnor2_4 c75 (.A(net11),
    .B(net819),
    .Y(net12));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(net395),
    .A1(net128),
    .A2(clknet_1_1__leaf_net354),
    .A3(clknet_1_1__leaf_net577),
    .S0(net748),
    .S1(net766),
    .X(net624));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net803),
    .A1(net482),
    .A2(net510),
    .A3(net788),
    .S0(net731),
    .S1(net760),
    .X(net625));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net575),
    .A1(net936),
    .A2(clknet_1_1__leaf_net142),
    .A3(net747),
    .S0(net765),
    .S1(net770),
    .X(net626));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net284),
    .A1(clknet_1_0__leaf_net560),
    .A2(net1008),
    .A3(clknet_1_1__leaf_net493),
    .S0(net787),
    .S1(clknet_1_1__leaf_net478),
    .X(net627));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net810),
    .A1(clknet_1_1__leaf_net376),
    .A2(net936),
    .A3(net818),
    .S0(net676),
    .S1(net771),
    .X(net628));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net19),
    .A1(net339),
    .A2(net334),
    .A3(net803),
    .S0(net679),
    .S1(net746),
    .X(net629));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net347),
    .A1(net69),
    .A2(net945),
    .A3(clknet_1_1__leaf_net695),
    .S0(net713),
    .S1(clknet_1_0__leaf_net735),
    .X(net630));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net787),
    .A1(net201),
    .A2(clknet_1_1__leaf_net120),
    .A3(net628),
    .S0(net621),
    .S1(net789),
    .X(net631));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net928),
    .A1(clknet_1_0__leaf_net577),
    .A2(net491),
    .A3(net631),
    .S0(clknet_1_1__leaf_net120),
    .S1(net769),
    .X(net632));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(clknet_1_1__leaf_net455),
    .A1(clknet_1_1__leaf_net103),
    .A2(net818),
    .A3(net519),
    .S0(net607),
    .S1(net803),
    .X(net633));
 sky130_fd_sc_hd__xnor2_4 c76 (.A(net7),
    .B(net5),
    .Y(net13));
 sky130_fd_sc_hd__mux4_2 c760 (.A0(net520),
    .A1(clknet_1_0__leaf_net268),
    .A2(net630),
    .A3(net704),
    .S0(net921),
    .S1(net740),
    .X(net634));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net295),
    .A1(net721),
    .A2(net754),
    .A3(net763),
    .S0(net767),
    .S1(net774));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net601),
    .A1(clknet_1_1__leaf_net478),
    .A2(net946),
    .A3(clknet_1_1__leaf_net515),
    .S0(clknet_1_1__leaf_net617),
    .S1(net773),
    .X(net635));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(net556),
    .A1(clknet_1_1__leaf_net548),
    .A2(net679),
    .A3(net680),
    .S0(net772),
    .S1(net775),
    .X(net636));
 sky130_fd_sc_hd__mux4_1 c764 (.A0(net629),
    .A1(net945),
    .A2(net195),
    .A3(net626),
    .S0(net636),
    .S1(net764));
 sky130_fd_sc_hd__xnor2_4 c77 (.A(net1011),
    .B(net1),
    .Y(net14));
 sky130_fd_sc_hd__xnor2_4 c78 (.A(net820),
    .B(net9),
    .Y(net15));
 sky130_fd_sc_hd__xnor2_4 c79 (.A(net15),
    .B(net12),
    .Y(net16));
 sky130_fd_sc_hd__a41o_4 c80 (.A1(net1),
    .A2(net16),
    .A3(net14),
    .A4(net791),
    .B1(net837),
    .X(net17));
 sky130_fd_sc_hd__a21bo_1 c81 (.A1(net14),
    .A2(net16),
    .B1_N(net824),
    .X(net18));
 sky130_fd_sc_hd__a41o_4 c82 (.A1(net16),
    .A2(net832),
    .A3(net13),
    .A4(net1),
    .B1(net795),
    .X(net860));
 sky130_fd_sc_hd__a41o_2 c83 (.A1(net18),
    .A2(net834),
    .A3(net916),
    .A4(net12),
    .B1(net802),
    .X(net19));
 sky130_fd_sc_hd__a31o_4 c84 (.A1(net904),
    .A2(net832),
    .A3(net4),
    .B1(net9),
    .X(net20));
 sky130_fd_sc_hd__xnor2_4 c85 (.A(net20),
    .B(net11),
    .Y(net872));
 sky130_fd_sc_hd__a31o_4 c86 (.A1(net872),
    .A2(net904),
    .A3(net10),
    .B1(net20),
    .X(net883));
 sky130_fd_sc_hd__xnor2_2 c87 (.A(net4),
    .B(net809),
    .Y(net21));
 sky130_fd_sc_hd__xnor2_4 c88 (.A(net788),
    .B(net883),
    .Y(net22));
 sky130_fd_sc_hd__xnor2_4 c89 (.A(net844),
    .B(net835),
    .Y(net23));
 sky130_fd_sc_hd__xnor2_4 c90 (.A(net796),
    .B(net14),
    .Y(net24));
 sky130_fd_sc_hd__xnor2_4 c91 (.A(net804),
    .B(net23),
    .Y(net25));
 sky130_fd_sc_hd__xnor2_4 c92 (.A(net22),
    .B(net25),
    .Y(net846));
 sky130_fd_sc_hd__xnor2_4 c93 (.A(net833),
    .B(net813),
    .Y(net845));
 sky130_fd_sc_hd__mux4_1 c94 (.A0(net792),
    .A1(net922),
    .A2(net16),
    .A3(net12),
    .S0(net13),
    .S1(net25),
    .X(net26));
 sky130_fd_sc_hd__xnor2_4 c95 (.A(net822),
    .B(net7),
    .Y(net27));
 sky130_fd_sc_hd__xnor2_2 c96 (.A(net24),
    .B(net10),
    .Y(net28));
 sky130_fd_sc_hd__xnor2_2 c97 (.A(net915),
    .B(net6),
    .Y(net29));
 sky130_fd_sc_hd__xnor2_2 c98 (.A(net915),
    .B(net6),
    .Y(net30));
 sky130_fd_sc_hd__xnor2_1 c99 (.A(net25),
    .B(net846),
    .Y(net31));
 sky130_fd_sc_hd__a41o_1 merge765 (.A1(net541),
    .A2(net527),
    .A3(net524),
    .A4(net531),
    .B1(net530),
    .X(net637));
 sky130_fd_sc_hd__mux4_1 merge766 (.A0(net21),
    .A1(clknet_1_0__leaf_net124),
    .A2(net911),
    .A3(net802),
    .S0(clknet_1_0__leaf_net127),
    .S1(net917),
    .X(net638));
 sky130_fd_sc_hd__mux4_1 merge767 (.A0(net808),
    .A1(net97),
    .A2(net215),
    .A3(net819),
    .S0(clknet_1_1__leaf_net125),
    .S1(net681),
    .X(net639));
 sky130_fd_sc_hd__buf_1 merge768 (.A(net780),
    .X(net640));
 sky130_fd_sc_hd__mux4_1 merge769 (.A0(net196),
    .A1(net189),
    .A2(net197),
    .A3(net203),
    .S0(net192),
    .S1(net190),
    .X(net641));
 sky130_fd_sc_hd__mux4_1 merge770 (.A0(net304),
    .A1(net346),
    .A2(net418),
    .A3(net445),
    .S0(net923),
    .S1(net211),
    .X(net642));
 sky130_fd_sc_hd__sdfbbn_1 merge771 (.CLK_N(clknet_4_0_0_clk),
    .D(net250),
    .RESET_B(net252),
    .SCE(net97),
    .SET_B(net714),
    .Q(net261),
    .Q_N(net643));
 sky130_fd_sc_hd__sdfbbp_1 merge772 (.CLK(clknet_4_2_0_clk),
    .D(net323),
    .RESET_B(net202),
    .SCD(clknet_1_0__leaf_net232),
    .SCE(clknet_1_0__leaf_net237),
    .SET_B(net853),
    .Q(net646),
    .Q_N(net645));
 sky130_fd_sc_hd__mux4_1 merge773 (.A0(clknet_1_1__leaf_net149),
    .A1(net918),
    .A2(net145),
    .A3(net157),
    .S0(net896),
    .S1(net150),
    .X(net647));
 sky130_fd_sc_hd__a41o_1 merge774 (.A1(net81),
    .A2(net97),
    .A3(clknet_1_0__leaf_net114),
    .A4(net111),
    .B1(net109),
    .X(net648));
 sky130_fd_sc_hd__a31o_1 merge775 (.A1(net791),
    .A2(net219),
    .A3(net933),
    .B1(net97),
    .X(net649));
 sky130_fd_sc_hd__a31o_1 merge776 (.A1(net797),
    .A2(net196),
    .A3(net791),
    .B1(net188),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_1 merge777 (.A(net699),
    .X(net651));
 sky130_fd_sc_hd__mux4_1 merge778 (.A0(net252),
    .A1(net929),
    .A2(net34),
    .A3(net15),
    .S0(net43),
    .S1(net969),
    .X(net652));
 sky130_fd_sc_hd__mux4_1 merge779 (.A0(net908),
    .A1(net159),
    .A2(clknet_1_0__leaf_net140),
    .A3(clknet_1_1__leaf_net132),
    .S0(clknet_1_0__leaf_net144),
    .S1(net674),
    .X(net653));
 sky130_fd_sc_hd__mux4_1 merge780 (.A0(clknet_1_0__leaf_net114),
    .A1(net106),
    .A2(net104),
    .A3(net207),
    .S0(clknet_1_0__leaf_net233),
    .S1(net930),
    .X(net654));
 sky130_fd_sc_hd__mux4_1 merge781 (.A0(net322),
    .A1(net808),
    .A2(net341),
    .A3(net327),
    .S0(net219),
    .S1(net691),
    .X(net655));
 sky130_fd_sc_hd__a41o_1 merge782 (.A1(net314),
    .A2(net418),
    .A3(net202),
    .A4(net185),
    .B1(net853),
    .X(net656));
 sky130_fd_sc_hd__mux4_1 merge783 (.A0(net235),
    .A1(net236),
    .A2(clknet_1_1__leaf_net237),
    .A3(net312),
    .S0(net302),
    .S1(net309),
    .X(net657));
 sky130_fd_sc_hd__mux4_1 merge784 (.A0(net526),
    .A1(net527),
    .A2(net524),
    .A3(clknet_1_0__leaf_net439),
    .S0(net787),
    .S1(clknet_1_0__leaf_net545),
    .X(net658));
 sky130_fd_sc_hd__mux4_1 merge785 (.A0(net74),
    .A1(net211),
    .A2(net301),
    .A3(net789),
    .S0(clknet_1_0__leaf_net233),
    .S1(net234),
    .X(net659));
 sky130_fd_sc_hd__mux4_2 merge786 (.A0(net843),
    .A1(clknet_1_1__leaf_net233),
    .A2(net869),
    .A3(net353),
    .S0(net997),
    .S1(net365),
    .X(net660));
 sky130_fd_sc_hd__mux4_1 merge787 (.A0(net175),
    .A1(net799),
    .A2(net172),
    .A3(net786),
    .S0(net42),
    .S1(net30),
    .X(net661));
 sky130_fd_sc_hd__mux4_1 merge788 (.A0(net349),
    .A1(net353),
    .A2(clknet_1_0__leaf_net354),
    .A3(net811),
    .S0(net201),
    .S1(net687),
    .X(net662));
 sky130_fd_sc_hd__mux4_1 merge789 (.A0(net304),
    .A1(net972),
    .A2(net894),
    .A3(net532),
    .S0(net71),
    .S1(net524),
    .X(net663));
 sky130_fd_sc_hd__mux4_1 merge790 (.A0(net535),
    .A1(net526),
    .A2(net527),
    .A3(net306),
    .S0(net536),
    .S1(net541),
    .X(net664));
 sky130_fd_sc_hd__dfrbp_1 merge791 (.CLK(clknet_4_11_0_clk),
    .D(net593),
    .RESET_B(net598),
    .Q(net666),
    .Q_N(net665));
 sky130_fd_sc_hd__dfrbp_1 merge792 (.CLK(clknet_4_0_0_clk),
    .D(net256),
    .RESET_B(net257),
    .Q(net668),
    .Q_N(net667));
 sky130_fd_sc_hd__dfrtn_1 merge793 (.CLK_N(clknet_4_8_0_clk),
    .D(net650),
    .RESET_B(net316),
    .Q(net669));
 sky130_fd_sc_hd__xnor2_1 merge794 (.A(net385),
    .B(net388),
    .Y(net670));
 sky130_fd_sc_hd__dfrtp_1 merge795 (.CLK(clknet_4_5_0_clk),
    .D(net55),
    .RESET_B(net61),
    .Q(net671));
 sky130_fd_sc_hd__dfrtp_1 merge796 (.CLK(clknet_4_12_0_clk),
    .D(net481),
    .Q(net492));
 sky130_fd_sc_hd__dfrtp_2 merge797 (.CLK(clknet_4_7_0_clk),
    .D(net397),
    .RESET_B(net399),
    .Q(net873));
 sky130_fd_sc_hd__xnor2_1 merge798 (.A(net648),
    .B(net654),
    .Y(net673));
 sky130_fd_sc_hd__dfsbp_1 merge799 (.CLK(clknet_4_4_0_clk),
    .D(net154),
    .SET_B(net160),
    .Q(net675),
    .Q_N(net674));
 sky130_fd_sc_hd__dfsbp_1 merge800 (.CLK(clknet_4_14_0_clk),
    .D(net602),
    .SET_B(net603),
    .Q(net677),
    .Q_N(net676));
 sky130_fd_sc_hd__dfstp_2 merge801 (.CLK(clknet_4_8_0_clk),
    .D(net430),
    .SET_B(net656),
    .Q(net678));
 sky130_fd_sc_hd__dfstp_1 merge802 (.CLK(clknet_4_15_0_clk),
    .D(net622),
    .SET_B(net623),
    .Q(net679));
 sky130_fd_sc_hd__dfstp_1 merge803 (.CLK(clknet_4_13_0_clk),
    .D(net501),
    .SET_B(net502),
    .Q(net680));
 sky130_fd_sc_hd__dlrbn_1 merge804 (.D(net297),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net298),
    .Q(net878),
    .Q_N(net879));
 sky130_fd_sc_hd__dlrbn_1 merge805 (.D(net226),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net225),
    .Q(net682),
    .Q_N(net681));
 sky130_fd_sc_hd__dlrbp_1 merge806 (.D(net466),
    .GATE(clknet_4_9_0_clk),
    .RESET_B(net473),
    .Q(net684),
    .Q_N(net683));
 sky130_fd_sc_hd__dlrbp_1 merge807 (.D(net637),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net658),
    .Q(net686),
    .Q_N(net685));
 sky130_fd_sc_hd__dlrtn_1 merge808 (.D(net359),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net364),
    .Q(net687));
 sky130_fd_sc_hd__dlrtn_1 merge809 (.D(net279),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net285),
    .Q(net688));
 sky130_fd_sc_hd__dlrtn_1 merge810 (.D(net169),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net171),
    .Q(net881));
 sky130_fd_sc_hd__dlrtp_1 merge811 (.D(net546),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net549),
    .Q(net689));
 sky130_fd_sc_hd__dlrtp_1 merge812 (.D(net133),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net638),
    .Q(net887));
 sky130_fd_sc_hd__dlrtp_1 merge813 (.D(net649),
    .GATE(clknet_4_2_0_clk),
    .RESET_B(net659),
    .Q(net690));
 sky130_fd_sc_hd__edfxbp_1 merge814 (.CLK(clknet_4_2_0_clk),
    .D(net212),
    .DE(net221),
    .Q(net692),
    .Q_N(net691));
 sky130_fd_sc_hd__edfxtp_1 merge815 (.CLK(clknet_4_1_0_clk),
    .D(net267),
    .DE(net299),
    .Q(net886));
 sky130_fd_sc_hd__sdlclkp_4 merge816 (.CLK(clknet_4_0_0_clk),
    .GATE(net99),
    .SCE(net673),
    .GCLK(net693));
 sky130_fd_sc_hd__sdlclkp_2 merge817 (.CLK(clknet_4_9_0_clk),
    .GATE(net476),
    .SCE(net479),
    .GCLK(net694));
 sky130_fd_sc_hd__sdlclkp_4 merge818 (.CLK(clknet_4_3_0_clk),
    .GATE(net670),
    .SCE(net620),
    .GCLK(net695));
 sky130_fd_sc_hd__dfrbp_1 merge819 (.CLK(clknet_4_7_0_clk),
    .D(net401),
    .RESET_B(net411),
    .Q(net697),
    .Q_N(net696));
 sky130_fd_sc_hd__dfrbp_1 merge820 (.CLK(clknet_4_10_0_clk),
    .D(net663),
    .RESET_B(net664),
    .Q(net699),
    .Q_N(net698));
 sky130_fd_sc_hd__dfrtn_1 merge821 (.CLK_N(clknet_4_12_0_clk),
    .D(net496),
    .RESET_B(net498),
    .Q(net700));
 sky130_fd_sc_hd__dfrtp_1 merge822 (.CLK(clknet_4_5_0_clk),
    .D(net165),
    .Q(net167));
 sky130_fd_sc_hd__dfrtp_4 merge823 (.CLK(clknet_4_1_0_clk),
    .D(net653),
    .RESET_B(net652),
    .Q(net702));
 sky130_fd_sc_hd__dfrtp_4 merge824 (.CLK(clknet_4_4_0_clk),
    .D(net647),
    .RESET_B(net138),
    .Q(net703));
 sky130_fd_sc_hd__dfsbp_1 merge825 (.CLK(clknet_4_7_0_clk),
    .D(net505),
    .SET_B(net506),
    .Q(net705),
    .Q_N(net704));
 sky130_fd_sc_hd__dfsbp_1 merge826 (.CLK(clknet_4_8_0_clk),
    .D(net641),
    .SET_B(net642),
    .Q(net707),
    .Q_N(net706));
 sky130_fd_sc_hd__dfstp_1 merge827 (.CLK(clknet_4_10_0_clk),
    .D(net558),
    .SET_B(net559),
    .Q(net708));
 sky130_fd_sc_hd__dfxbp_1 s828 (.CLK(clknet_4_5_0_clk),
    .D(net164),
    .Q(net710),
    .Q_N(net709));
 sky130_fd_sc_hd__dfxbp_1 s829 (.CLK(clknet_4_5_0_clk),
    .D(net173),
    .Q(net712),
    .Q_N(net711));
 sky130_fd_sc_hd__dfxtp_1 s830 (.CLK(clknet_4_5_0_clk),
    .D(net181),
    .Q(net859));
 sky130_fd_sc_hd__dfxtp_4 s831 (.CLK(clknet_4_2_0_clk),
    .D(net216),
    .Q(net713));
 sky130_fd_sc_hd__dfxtp_2 s832 (.CLK(clknet_4_0_0_clk),
    .D(net229),
    .Q(net714));
 sky130_fd_sc_hd__dlclkp_1 s833 (.CLK(clknet_4_0_0_clk),
    .GATE(net240),
    .GCLK(net715));
 sky130_fd_sc_hd__dlclkp_2 s834 (.CLK(clknet_4_3_0_clk),
    .GATE(net246),
    .GCLK(net716));
 sky130_fd_sc_hd__dlclkp_4 s835 (.CLK(clknet_4_5_0_clk),
    .GATE(net286),
    .GCLK(net863));
 sky130_fd_sc_hd__dlxbn_1 s836 (.D(net293),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net718),
    .Q_N(net717));
 sky130_fd_sc_hd__dlxbn_1 s837 (.D(net296),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net875),
    .Q_N(net719));
 sky130_fd_sc_hd__dlxbp_1 s838 (.D(net363),
    .GATE(clknet_4_14_0_clk),
    .Q(net721),
    .Q_N(net720));
 sky130_fd_sc_hd__dlxtn_1 s839 (.D(net370),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net722));
 sky130_fd_sc_hd__dlxtn_1 s840 (.D(net375),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net723));
 sky130_fd_sc_hd__dlxtn_1 s841 (.D(net381),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net724));
 sky130_fd_sc_hd__dlxtp_1 s842 (.D(net394),
    .GATE(clknet_4_6_0_clk),
    .Q(net725));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s843 (.D(net398),
    .SLEEP_B(clknet_4_6_0_clk),
    .Q(net726));
 sky130_fd_sc_hd__dfxbp_1 s844 (.CLK(clknet_4_7_0_clk),
    .D(net400),
    .Q(net728),
    .Q_N(net727));
 sky130_fd_sc_hd__dfxbp_1 s845 (.CLK(clknet_4_7_0_clk),
    .D(net404),
    .Q(net729));
 sky130_fd_sc_hd__dfxtp_1 s846 (.CLK(clknet_4_7_0_clk),
    .D(net407),
    .Q(net730));
 sky130_fd_sc_hd__dfxtp_2 s847 (.CLK(clknet_4_7_0_clk),
    .D(net409),
    .Q(net731));
 sky130_fd_sc_hd__dfxtp_1 s848 (.CLK(clknet_4_7_0_clk),
    .D(net410),
    .Q(net732));
 sky130_fd_sc_hd__dlclkp_1 s849 (.CLK(clknet_4_8_0_clk),
    .GATE(net434),
    .GCLK(net733));
 sky130_fd_sc_hd__dlclkp_2 s850 (.CLK(clknet_4_9_0_clk),
    .GATE(net467),
    .GCLK(net734));
 sky130_fd_sc_hd__dlclkp_4 s851 (.CLK(clknet_4_12_0_clk),
    .GATE(net490),
    .GCLK(net735));
 sky130_fd_sc_hd__dlxbn_1 s852 (.D(net497),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net737),
    .Q_N(net736));
 sky130_fd_sc_hd__dlxbn_1 s853 (.D(net499),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net854),
    .Q_N(net738));
 sky130_fd_sc_hd__dlxbp_1 s854 (.D(net507),
    .GATE(clknet_4_12_0_clk),
    .Q(net739));
 sky130_fd_sc_hd__dlxtn_1 s855 (.D(net508),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net740));
 sky130_fd_sc_hd__dlxtn_1 s856 (.D(net509),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net741));
 sky130_fd_sc_hd__dlxtn_1 s857 (.D(net511),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net742));
 sky130_fd_sc_hd__dlxtp_1 s858 (.D(net512),
    .GATE(clknet_4_13_0_clk),
    .Q(net743));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s859 (.D(net513),
    .SLEEP_B(clknet_4_13_0_clk),
    .Q(net744));
 sky130_fd_sc_hd__dfxbp_1 s860 (.CLK(clknet_4_13_0_clk),
    .D(net517),
    .Q(net745));
 sky130_fd_sc_hd__dfxbp_1 s861 (.CLK(clknet_4_13_0_clk),
    .D(net518),
    .Q(net746));
 sky130_fd_sc_hd__dfxtp_1 s862 (.CLK(clknet_4_13_0_clk),
    .D(net521),
    .Q(net747));
 sky130_fd_sc_hd__dfxtp_1 s863 (.CLK(clknet_4_13_0_clk),
    .D(net522),
    .Q(net748));
 sky130_fd_sc_hd__dfxtp_1 s864 (.CLK(clknet_4_10_0_clk),
    .D(net568),
    .Q(net749));
 sky130_fd_sc_hd__dlclkp_1 s865 (.CLK(clknet_4_11_0_clk),
    .GATE(net569),
    .GCLK(net750));
 sky130_fd_sc_hd__dlclkp_2 s866 (.CLK(clknet_4_11_0_clk),
    .GATE(net573),
    .GCLK(net751));
 sky130_fd_sc_hd__dlclkp_4 s867 (.CLK(clknet_4_14_0_clk),
    .GATE(net576),
    .GCLK(net752));
 sky130_fd_sc_hd__dlxbn_1 s868 (.D(net588),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net754),
    .Q_N(net753));
 sky130_fd_sc_hd__dlxbn_1 s869 (.D(net591),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net756),
    .Q_N(net755));
 sky130_fd_sc_hd__dlxbp_1 s870 (.D(net594),
    .GATE(clknet_4_11_0_clk),
    .Q(net758),
    .Q_N(net757));
 sky130_fd_sc_hd__dlxtn_1 s871 (.D(net599),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net759));
 sky130_fd_sc_hd__dlxtn_1 s872 (.D(net604),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net760));
 sky130_fd_sc_hd__dlxtn_1 s873 (.D(net605),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net761));
 sky130_fd_sc_hd__dlxtp_1 s874 (.D(net608),
    .GATE(clknet_4_15_0_clk),
    .Q(net762));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s875 (.D(net609),
    .SLEEP_B(clknet_4_14_0_clk),
    .Q(net763));
 sky130_fd_sc_hd__dfxbp_1 s876 (.CLK(clknet_4_13_0_clk),
    .D(net611),
    .Q(net764));
 sky130_fd_sc_hd__dfxbp_1 s877 (.CLK(clknet_4_15_0_clk),
    .D(net613),
    .Q(net765));
 sky130_fd_sc_hd__dfxtp_1 s878 (.CLK(clknet_4_13_0_clk),
    .D(net614),
    .Q(net766));
 sky130_fd_sc_hd__dfxtp_1 s879 (.CLK(clknet_4_14_0_clk),
    .D(net615),
    .Q(net767));
 sky130_fd_sc_hd__dfxtp_1 s880 (.CLK(clknet_4_15_0_clk),
    .D(net616),
    .Q(net768));
 sky130_fd_sc_hd__dlclkp_1 s881 (.CLK(clknet_4_13_0_clk),
    .GATE(net624),
    .GCLK(net769));
 sky130_fd_sc_hd__dlclkp_2 s882 (.CLK(clknet_4_13_0_clk),
    .GATE(net625),
    .GCLK(net770));
 sky130_fd_sc_hd__dlclkp_4 s883 (.CLK(clknet_4_12_0_clk),
    .GATE(net627),
    .GCLK(net771));
 sky130_fd_sc_hd__dlxbn_1 s884 (.D(net632),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net772));
 sky130_fd_sc_hd__dlxbn_1 s885 (.D(net633),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net773));
 sky130_fd_sc_hd__dlxbp_1 s886 (.D(net634),
    .GATE(clknet_4_15_0_clk),
    .Q(net774));
 sky130_fd_sc_hd__dlxtn_1 s887 (.D(net635),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net775));
 sky130_fd_sc_hd__dlxtn_1 s888 (.D(net639),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net776));
 sky130_fd_sc_hd__dlxtn_1 s889 (.D(net655),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net777));
 sky130_fd_sc_hd__dlxtp_1 s890 (.D(net657),
    .GATE(clknet_4_2_0_clk),
    .Q(net778));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s891 (.D(net660),
    .SLEEP_B(clknet_4_3_0_clk),
    .Q(net779));
 sky130_fd_sc_hd__dfxbp_1 s892 (.CLK(clknet_4_5_0_clk),
    .D(net661),
    .Q(net781),
    .Q_N(net780));
 sky130_fd_sc_hd__dfxbp_1 s893 (.CLK(clknet_4_9_0_clk),
    .D(net662),
    .Q(net783),
    .Q_N(net782));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_12 input1 (.A(in0),
    .X(net644));
 sky130_fd_sc_hd__buf_2 input2 (.A(in1),
    .X(net784));
 sky130_fd_sc_hd__buf_8 input3 (.A(in10),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(in11),
    .X(net786));
 sky130_fd_sc_hd__buf_4 input5 (.A(in12),
    .X(net787));
 sky130_fd_sc_hd__buf_4 input6 (.A(in13),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_8 input7 (.A(in14),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_8 input8 (.A(in15),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_8 input9 (.A(in16),
    .X(net791));
 sky130_fd_sc_hd__buf_8 input10 (.A(in17),
    .X(net792));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(in18),
    .X(net793));
 sky130_fd_sc_hd__clkbuf_8 input12 (.A(in19),
    .X(net794));
 sky130_fd_sc_hd__buf_6 input13 (.A(in2),
    .X(net795));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(in20),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(in21),
    .X(net797));
 sky130_fd_sc_hd__buf_4 input16 (.A(in22),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_8 input17 (.A(in23),
    .X(net799));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(in24),
    .X(net800));
 sky130_fd_sc_hd__buf_4 input19 (.A(in25),
    .X(net801));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(in26),
    .X(net802));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(in27),
    .X(net803));
 sky130_fd_sc_hd__buf_6 input22 (.A(in28),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(in29),
    .X(net805));
 sky130_fd_sc_hd__buf_4 input24 (.A(in3),
    .X(net806));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(in30),
    .X(net807));
 sky130_fd_sc_hd__buf_2 input26 (.A(in31),
    .X(net808));
 sky130_fd_sc_hd__clkbuf_4 input27 (.A(in32),
    .X(net809));
 sky130_fd_sc_hd__buf_4 input28 (.A(in33),
    .X(net810));
 sky130_fd_sc_hd__buf_2 input29 (.A(in34),
    .X(net811));
 sky130_fd_sc_hd__buf_2 input30 (.A(in35),
    .X(net812));
 sky130_fd_sc_hd__buf_8 input31 (.A(in36),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(in37),
    .X(net814));
 sky130_fd_sc_hd__buf_4 input33 (.A(in38),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(in39),
    .X(net816));
 sky130_fd_sc_hd__buf_12 input35 (.A(in4),
    .X(net817));
 sky130_fd_sc_hd__buf_6 input36 (.A(in40),
    .X(net818));
 sky130_fd_sc_hd__buf_4 input37 (.A(in41),
    .X(net819));
 sky130_fd_sc_hd__clkbuf_8 input38 (.A(in42),
    .X(net820));
 sky130_fd_sc_hd__clkbuf_4 input39 (.A(in43),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_4 input40 (.A(in44),
    .X(net822));
 sky130_fd_sc_hd__buf_2 input41 (.A(in45),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(in46),
    .X(net824));
 sky130_fd_sc_hd__buf_2 input43 (.A(in47),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(in48),
    .X(net826));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(in49),
    .X(net827));
 sky130_fd_sc_hd__clkbuf_8 input46 (.A(in5),
    .X(net828));
 sky130_fd_sc_hd__clkbuf_8 input47 (.A(in50),
    .X(net829));
 sky130_fd_sc_hd__buf_1 input48 (.A(in51),
    .X(net830));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(in52),
    .X(net831));
 sky130_fd_sc_hd__buf_4 input50 (.A(in53),
    .X(net832));
 sky130_fd_sc_hd__buf_2 input51 (.A(in54),
    .X(net833));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(in55),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(in56),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(in57),
    .X(net836));
 sky130_fd_sc_hd__buf_2 input55 (.A(in58),
    .X(net837));
 sky130_fd_sc_hd__buf_2 input56 (.A(in59),
    .X(net838));
 sky130_fd_sc_hd__buf_6 input57 (.A(in6),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_4 input58 (.A(in60),
    .X(net840));
 sky130_fd_sc_hd__clkbuf_4 input59 (.A(net1012),
    .X(net841));
 sky130_fd_sc_hd__buf_4 input60 (.A(in7),
    .X(net842));
 sky130_fd_sc_hd__buf_4 input61 (.A(in8),
    .X(net843));
 sky130_fd_sc_hd__clkbuf_8 input62 (.A(in9),
    .X(net844));
 sky130_fd_sc_hd__buf_2 output63 (.A(net922),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output64 (.A(net846),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output65 (.A(net847),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output66 (.A(net848),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output67 (.A(net849),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output68 (.A(net850),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output69 (.A(net851),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output70 (.A(net852),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output71 (.A(net853),
    .X(out2));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net854),
    .X(out20));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net855),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output74 (.A(net856),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output75 (.A(net857),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output76 (.A(net858),
    .X(out25));
 sky130_fd_sc_hd__buf_2 output77 (.A(net859),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output78 (.A(net860),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output79 (.A(net861),
    .X(out29));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net862),
    .X(out3));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(clknet_1_1__leaf_net863),
    .X(out30));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net864),
    .X(out31));
 sky130_fd_sc_hd__buf_2 output83 (.A(net865),
    .X(out32));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(clknet_1_1__leaf_net866),
    .X(out33));
 sky130_fd_sc_hd__buf_2 output85 (.A(net867),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output86 (.A(net868),
    .X(out36));
 sky130_fd_sc_hd__buf_2 output87 (.A(net869),
    .X(out37));
 sky130_fd_sc_hd__buf_2 output88 (.A(net870),
    .X(out38));
 sky130_fd_sc_hd__buf_2 output89 (.A(net871),
    .X(out41));
 sky130_fd_sc_hd__buf_2 output90 (.A(net872),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output91 (.A(net873),
    .X(out43));
 sky130_fd_sc_hd__buf_2 output92 (.A(net874),
    .X(out44));
 sky130_fd_sc_hd__buf_2 output93 (.A(net875),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output94 (.A(net876),
    .X(out46));
 sky130_fd_sc_hd__buf_2 output95 (.A(net877),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output96 (.A(net878),
    .X(out48));
 sky130_fd_sc_hd__buf_2 output97 (.A(net879),
    .X(out49));
 sky130_fd_sc_hd__buf_2 output98 (.A(net880),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output99 (.A(net881),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output100 (.A(net882),
    .X(out51));
 sky130_fd_sc_hd__buf_2 output101 (.A(net883),
    .X(out52));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(clknet_1_0__leaf_net884),
    .X(out53));
 sky130_fd_sc_hd__buf_2 output103 (.A(net885),
    .X(out54));
 sky130_fd_sc_hd__buf_2 output104 (.A(net886),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output105 (.A(net887),
    .X(out56));
 sky130_fd_sc_hd__buf_2 output106 (.A(net888),
    .X(out57));
 sky130_fd_sc_hd__buf_2 output107 (.A(net889),
    .X(out59));
 sky130_fd_sc_hd__clkbuf_1 output108 (.A(clknet_1_1__leaf_net890),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output109 (.A(net891),
    .X(out60));
 sky130_fd_sc_hd__buf_2 output110 (.A(net892),
    .X(out61));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(net893),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_4 output112 (.A(net894),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_4 fanout113 (.A(net563),
    .X(net895));
 sky130_fd_sc_hd__clkbuf_4 fanout114 (.A(net856),
    .X(net896));
 sky130_fd_sc_hd__buf_4 max_cap115 (.A(net874),
    .X(net897));
 sky130_fd_sc_hd__buf_6 fanout116 (.A(net195),
    .X(net898));
 sky130_fd_sc_hd__buf_4 max_cap117 (.A(net308),
    .X(net899));
 sky130_fd_sc_hd__clkbuf_8 fanout118 (.A(net191),
    .X(net900));
 sky130_fd_sc_hd__buf_4 max_cap119 (.A(net206),
    .X(net901));
 sky130_fd_sc_hd__buf_12 fanout120 (.A(net80),
    .X(net902));
 sky130_fd_sc_hd__buf_4 max_cap121 (.A(net186),
    .X(net903));
 sky130_fd_sc_hd__buf_4 fanout122 (.A(net19),
    .X(net904));
 sky130_fd_sc_hd__buf_12 fanout123 (.A(net71),
    .X(net905));
 sky130_fd_sc_hd__buf_6 fanout124 (.A(net961),
    .X(net906));
 sky130_fd_sc_hd__buf_12 max_cap125 (.A(net70),
    .X(net907));
 sky130_fd_sc_hd__buf_4 max_cap126 (.A(net83),
    .X(net908));
 sky130_fd_sc_hd__buf_6 fanout127 (.A(net910),
    .X(net909));
 sky130_fd_sc_hd__buf_8 fanout128 (.A(net912),
    .X(net910));
 sky130_fd_sc_hd__buf_4 fanout129 (.A(net912),
    .X(net911));
 sky130_fd_sc_hd__buf_6 fanout130 (.A(net72),
    .X(net912));
 sky130_fd_sc_hd__buf_4 max_cap131 (.A(net914),
    .X(net913));
 sky130_fd_sc_hd__buf_8 max_cap132 (.A(net68),
    .X(net914));
 sky130_fd_sc_hd__buf_4 max_cap133 (.A(net27),
    .X(net915));
 sky130_fd_sc_hd__buf_4 max_cap134 (.A(net5),
    .X(net916));
 sky130_fd_sc_hd__clkbuf_4 fanout135 (.A(net918),
    .X(net917));
 sky130_fd_sc_hd__buf_4 fanout136 (.A(net128),
    .X(net918));
 sky130_fd_sc_hd__buf_4 max_cap137 (.A(net69),
    .X(net919));
 sky130_fd_sc_hd__buf_8 max_cap138 (.A(net65),
    .X(net920));
 sky130_fd_sc_hd__clkbuf_4 fanout139 (.A(net724),
    .X(net921));
 sky130_fd_sc_hd__clkbuf_4 fanout140 (.A(net845),
    .X(net922));
 sky130_fd_sc_hd__clkbuf_4 fanout141 (.A(net967),
    .X(net923));
 sky130_fd_sc_hd__buf_4 fanout142 (.A(net339),
    .X(net924));
 sky130_fd_sc_hd__buf_4 max_cap143 (.A(net877),
    .X(net925));
 sky130_fd_sc_hd__buf_4 max_cap144 (.A(net64),
    .X(net926));
 sky130_fd_sc_hd__buf_4 wire145 (.A(net63),
    .X(net927));
 sky130_fd_sc_hd__buf_4 fanout146 (.A(net62),
    .X(net928));
 sky130_fd_sc_hd__buf_4 fanout147 (.A(net836),
    .X(net929));
 sky130_fd_sc_hd__buf_6 fanout148 (.A(net1008),
    .X(net930));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(net950),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(net950),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(net950),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(net950),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(net950),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(net948),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(net949),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(net948),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(net948),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net752 (.A(net752),
    .X(clknet_0_net752));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net752 (.A(clknet_0_net752),
    .X(clknet_1_0__leaf_net752));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net752 (.A(clknet_0_net752),
    .X(clknet_1_1__leaf_net752));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net751 (.A(net751),
    .X(clknet_0_net751));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net751 (.A(clknet_0_net751),
    .X(clknet_1_0__leaf_net751));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net751 (.A(clknet_0_net751),
    .X(clknet_1_1__leaf_net751));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net596 (.A(net596),
    .X(clknet_0_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net596 (.A(clknet_0_net596),
    .X(clknet_1_0__leaf_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net596 (.A(clknet_0_net596),
    .X(clknet_1_1__leaf_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net750 (.A(net750),
    .X(clknet_0_net750));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net750 (.A(clknet_0_net750),
    .X(clknet_1_0__leaf_net750));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net750 (.A(clknet_0_net750),
    .X(clknet_1_1__leaf_net750));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net617 (.A(net617),
    .X(clknet_0_net617));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net617 (.A(clknet_0_net617),
    .X(clknet_1_0__leaf_net617));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net617 (.A(clknet_0_net617),
    .X(clknet_1_1__leaf_net617));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net695 (.A(net695),
    .X(clknet_0_net695));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net695 (.A(clknet_0_net695),
    .X(clknet_1_0__leaf_net695));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net695 (.A(clknet_0_net695),
    .X(clknet_1_1__leaf_net695));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net735 (.A(net735),
    .X(clknet_0_net735));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net735 (.A(clknet_0_net735),
    .X(clknet_1_0__leaf_net735));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net735 (.A(clknet_0_net735),
    .X(clknet_1_1__leaf_net735));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net734 (.A(net734),
    .X(clknet_0_net734));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net734 (.A(clknet_0_net734),
    .X(clknet_1_0__leaf_net734));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net734 (.A(clknet_0_net734),
    .X(clknet_1_1__leaf_net734));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net694 (.A(net694),
    .X(clknet_0_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net694 (.A(clknet_0_net694),
    .X(clknet_1_0__leaf_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net694 (.A(clknet_0_net694),
    .X(clknet_1_1__leaf_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net582 (.A(net582),
    .X(clknet_0_net582));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net582 (.A(clknet_0_net582),
    .X(clknet_1_0__leaf_net582));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net582 (.A(clknet_0_net582),
    .X(clknet_1_1__leaf_net582));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net471 (.A(net471),
    .X(clknet_0_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net471 (.A(clknet_0_net471),
    .X(clknet_1_0__leaf_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net471 (.A(clknet_0_net471),
    .X(clknet_1_1__leaf_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net472 (.A(net472),
    .X(clknet_0_net472));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net472 (.A(clknet_0_net472),
    .X(clknet_1_0__leaf_net472));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net472 (.A(clknet_0_net472),
    .X(clknet_1_1__leaf_net472));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net733 (.A(net733),
    .X(clknet_0_net733));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net733 (.A(clknet_0_net733),
    .X(clknet_1_0__leaf_net733));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net733 (.A(clknet_0_net733),
    .X(clknet_1_1__leaf_net733));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net448 (.A(net448),
    .X(clknet_0_net448));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net448 (.A(clknet_0_net448),
    .X(clknet_1_0__leaf_net448));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net448 (.A(clknet_0_net448),
    .X(clknet_1_1__leaf_net448));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net485 (.A(net485),
    .X(clknet_0_net485));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net485 (.A(clknet_0_net485),
    .X(clknet_1_0__leaf_net485));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net485 (.A(clknet_0_net485),
    .X(clknet_1_1__leaf_net485));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net438 (.A(net438),
    .X(clknet_0_net438));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net438 (.A(clknet_0_net438),
    .X(clknet_1_0__leaf_net438));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net438 (.A(clknet_0_net438),
    .X(clknet_1_1__leaf_net438));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net577 (.A(net577),
    .X(clknet_0_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net577 (.A(clknet_0_net577),
    .X(clknet_1_0__leaf_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net577 (.A(clknet_0_net577),
    .X(clknet_1_1__leaf_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net548 (.A(net548),
    .X(clknet_0_net548));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net548 (.A(clknet_0_net548),
    .X(clknet_1_0__leaf_net548));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net548 (.A(clknet_0_net548),
    .X(clknet_1_1__leaf_net548));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net437 (.A(net437),
    .X(clknet_0_net437));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net437 (.A(clknet_0_net437),
    .X(clknet_1_0__leaf_net437));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net437 (.A(clknet_0_net437),
    .X(clknet_1_1__leaf_net437));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net455 (.A(net455),
    .X(clknet_0_net455));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net455 (.A(clknet_0_net455),
    .X(clknet_1_0__leaf_net455));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net455 (.A(clknet_0_net455),
    .X(clknet_1_1__leaf_net455));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net478 (.A(net478),
    .X(clknet_0_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net478 (.A(clknet_0_net478),
    .X(clknet_1_0__leaf_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net478 (.A(clknet_0_net478),
    .X(clknet_1_1__leaf_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net443 (.A(net443),
    .X(clknet_0_net443));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net443 (.A(clknet_0_net443),
    .X(clknet_1_0__leaf_net443));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net443 (.A(clknet_0_net443),
    .X(clknet_1_1__leaf_net443));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net439 (.A(net439),
    .X(clknet_0_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net439 (.A(clknet_0_net439),
    .X(clknet_1_0__leaf_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net439 (.A(clknet_0_net439),
    .X(clknet_1_1__leaf_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net545 (.A(net545),
    .X(clknet_0_net545));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net545 (.A(clknet_0_net545),
    .X(clknet_1_0__leaf_net545));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net545 (.A(clknet_0_net545),
    .X(clknet_1_1__leaf_net545));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net440 (.A(net440),
    .X(clknet_0_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net440 (.A(clknet_0_net440),
    .X(clknet_1_0__leaf_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net440 (.A(clknet_0_net440),
    .X(clknet_1_1__leaf_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net863 (.A(net863),
    .X(clknet_0_net863));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net863 (.A(clknet_0_net863),
    .X(clknet_1_0__leaf_net863));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net863 (.A(clknet_0_net863),
    .X(clknet_1_1__leaf_net863));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net292 (.A(net292),
    .X(clknet_0_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net292 (.A(clknet_0_net292),
    .X(clknet_1_0__leaf_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net292 (.A(clknet_0_net292),
    .X(clknet_1_1__leaf_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net290 (.A(net290),
    .X(clknet_0_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net290 (.A(clknet_0_net290),
    .X(clknet_1_0__leaf_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net290 (.A(clknet_0_net290),
    .X(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net716 (.A(net716),
    .X(clknet_0_net716));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net716 (.A(clknet_0_net716),
    .X(clknet_1_0__leaf_net716));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net716 (.A(clknet_0_net716),
    .X(clknet_1_1__leaf_net716));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net249 (.A(net249),
    .X(clknet_0_net249));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net249 (.A(clknet_0_net249),
    .X(clknet_1_0__leaf_net249));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net249 (.A(clknet_0_net249),
    .X(clknet_1_1__leaf_net249));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net266 (.A(net266),
    .X(clknet_0_net266));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net266 (.A(clknet_0_net266),
    .X(clknet_1_0__leaf_net266));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net266 (.A(clknet_0_net266),
    .X(clknet_1_1__leaf_net266));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net270 (.A(net270),
    .X(clknet_0_net270));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net270 (.A(clknet_0_net270),
    .X(clknet_1_0__leaf_net270));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net270 (.A(clknet_0_net270),
    .X(clknet_1_1__leaf_net270));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net387 (.A(net387),
    .X(clknet_0_net387));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net387 (.A(clknet_0_net387),
    .X(clknet_1_0__leaf_net387));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net387 (.A(clknet_0_net387),
    .X(clknet_1_1__leaf_net387));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net269 (.A(net269),
    .X(clknet_0_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net269 (.A(clknet_0_net269),
    .X(clknet_1_0__leaf_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net269 (.A(clknet_0_net269),
    .X(clknet_1_1__leaf_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net715 (.A(net715),
    .X(clknet_0_net715));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net715 (.A(clknet_0_net715),
    .X(clknet_1_0__leaf_net715));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net715 (.A(clknet_0_net715),
    .X(clknet_1_1__leaf_net715));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net251 (.A(net251),
    .X(clknet_0_net251));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net251 (.A(clknet_0_net251),
    .X(clknet_1_0__leaf_net251));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net251 (.A(clknet_0_net251),
    .X(clknet_1_1__leaf_net251));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net693 (.A(net693),
    .X(clknet_0_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net693 (.A(clknet_0_net693),
    .X(clknet_1_0__leaf_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net693 (.A(clknet_0_net693),
    .X(clknet_1_1__leaf_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net237 (.A(net237),
    .X(clknet_0_net237));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net237 (.A(clknet_0_net237),
    .X(clknet_1_0__leaf_net237));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net237 (.A(clknet_0_net237),
    .X(clknet_1_1__leaf_net237));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net241 (.A(net241),
    .X(clknet_0_net241));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net241 (.A(clknet_0_net241),
    .X(clknet_1_0__leaf_net241));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net241 (.A(clknet_0_net241),
    .X(clknet_1_1__leaf_net241));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net121 (.A(net121),
    .X(clknet_0_net121));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net121 (.A(clknet_0_net121),
    .X(clknet_1_0__leaf_net121));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net121 (.A(clknet_0_net121),
    .X(clknet_1_1__leaf_net121));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net230 (.A(net230),
    .X(clknet_0_net230));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net230 (.A(clknet_0_net230),
    .X(clknet_1_0__leaf_net230));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net230 (.A(clknet_0_net230),
    .X(clknet_1_1__leaf_net230));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net357 (.A(net357),
    .X(clknet_0_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net357 (.A(clknet_0_net357),
    .X(clknet_1_0__leaf_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net357 (.A(clknet_0_net357),
    .X(clknet_1_1__leaf_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net360 (.A(net360),
    .X(clknet_0_net360));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net360 (.A(clknet_0_net360),
    .X(clknet_1_0__leaf_net360));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net360 (.A(clknet_0_net360),
    .X(clknet_1_1__leaf_net360));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net366 (.A(net366),
    .X(clknet_0_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net366 (.A(clknet_0_net366),
    .X(clknet_1_0__leaf_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net366 (.A(clknet_0_net366),
    .X(clknet_1_1__leaf_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net232 (.A(net232),
    .X(clknet_0_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net232 (.A(clknet_0_net232),
    .X(clknet_1_0__leaf_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net232 (.A(clknet_0_net232),
    .X(clknet_1_1__leaf_net232));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net890 (.A(net890),
    .X(clknet_0_net890));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net890 (.A(clknet_0_net890),
    .X(clknet_1_0__leaf_net890));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net890 (.A(clknet_0_net890),
    .X(clknet_1_1__leaf_net890));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net233 (.A(net233),
    .X(clknet_0_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net233 (.A(clknet_0_net233),
    .X(clknet_1_0__leaf_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net233 (.A(clknet_0_net233),
    .X(clknet_1_1__leaf_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net117 (.A(net117),
    .X(clknet_0_net117));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net117 (.A(clknet_0_net117),
    .X(clknet_1_0__leaf_net117));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net117 (.A(clknet_0_net117),
    .X(clknet_1_1__leaf_net117));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net469 (.A(net469),
    .X(clknet_0_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net469 (.A(clknet_0_net469),
    .X(clknet_1_0__leaf_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net469 (.A(clknet_0_net469),
    .X(clknet_1_1__leaf_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net124 (.A(net124),
    .X(clknet_0_net124));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net124 (.A(clknet_0_net124),
    .X(clknet_1_0__leaf_net124));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net124 (.A(clknet_0_net124),
    .X(clknet_1_1__leaf_net124));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net118 (.A(net118),
    .X(clknet_0_net118));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net118 (.A(clknet_0_net118),
    .X(clknet_1_0__leaf_net118));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net118 (.A(clknet_0_net118),
    .X(clknet_1_1__leaf_net118));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net132 (.A(net132),
    .X(clknet_0_net132));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net132 (.A(clknet_0_net132),
    .X(clknet_1_0__leaf_net132));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net132 (.A(clknet_0_net132),
    .X(clknet_1_1__leaf_net132));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net140 (.A(net140),
    .X(clknet_0_net140));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net140 (.A(clknet_0_net140),
    .X(clknet_1_0__leaf_net140));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net140 (.A(clknet_0_net140),
    .X(clknet_1_1__leaf_net140));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net866 (.A(net866),
    .X(clknet_0_net866));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net866 (.A(clknet_0_net866),
    .X(clknet_1_0__leaf_net866));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net866 (.A(clknet_0_net866),
    .X(clknet_1_1__leaf_net866));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net412 (.A(net412),
    .X(clknet_0_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net412 (.A(clknet_0_net412),
    .X(clknet_1_0__leaf_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net412 (.A(clknet_0_net412),
    .X(clknet_1_1__leaf_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net144 (.A(net144),
    .X(clknet_0_net144));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net144 (.A(clknet_0_net144),
    .X(clknet_1_0__leaf_net144));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net144 (.A(clknet_0_net144),
    .X(clknet_1_1__leaf_net144));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net143 (.A(net143),
    .X(clknet_0_net143));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net143 (.A(clknet_0_net143),
    .X(clknet_1_0__leaf_net143));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net143 (.A(clknet_0_net143),
    .X(clknet_1_1__leaf_net143));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net142 (.A(net142),
    .X(clknet_0_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net142 (.A(clknet_0_net142),
    .X(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net142 (.A(clknet_0_net142),
    .X(clknet_1_1__leaf_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net493 (.A(net493),
    .X(clknet_0_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net493 (.A(clknet_0_net493),
    .X(clknet_1_0__leaf_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net493 (.A(clknet_0_net493),
    .X(clknet_1_1__leaf_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net282 (.A(net282),
    .X(clknet_0_net282));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net282 (.A(clknet_0_net282),
    .X(clknet_1_0__leaf_net282));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net282 (.A(clknet_0_net282),
    .X(clknet_1_1__leaf_net282));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net149 (.A(net149),
    .X(clknet_0_net149));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net149 (.A(clknet_0_net149),
    .X(clknet_1_0__leaf_net149));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net149 (.A(clknet_0_net149),
    .X(clknet_1_1__leaf_net149));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net134 (.A(net134),
    .X(clknet_0_net134));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net134 (.A(clknet_0_net134),
    .X(clknet_1_0__leaf_net134));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net134 (.A(clknet_0_net134),
    .X(clknet_1_1__leaf_net134));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net137 (.A(net137),
    .X(clknet_0_net137));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net137 (.A(clknet_0_net137),
    .X(clknet_1_0__leaf_net137));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net137 (.A(net958),
    .X(clknet_1_1__leaf_net137));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net263 (.A(net263),
    .X(clknet_0_net263));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net263 (.A(clknet_0_net263),
    .X(clknet_1_0__leaf_net263));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net263 (.A(net957),
    .X(clknet_1_1__leaf_net263));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net268 (.A(net268),
    .X(clknet_0_net268));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net268 (.A(clknet_0_net268),
    .X(clknet_1_0__leaf_net268));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net268 (.A(net953),
    .X(clknet_1_1__leaf_net268));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net489 (.A(net489),
    .X(clknet_0_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_0__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_1__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net383 (.A(net383),
    .X(clknet_0_net383));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net383 (.A(clknet_0_net383),
    .X(clknet_1_0__leaf_net383));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net383 (.A(clknet_0_net383),
    .X(clknet_1_1__leaf_net383));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net386 (.A(net386),
    .X(clknet_0_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net386 (.A(clknet_0_net386),
    .X(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net386 (.A(clknet_0_net386),
    .X(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net382 (.A(net382),
    .X(clknet_0_net382));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net382 (.A(clknet_0_net382),
    .X(clknet_1_0__leaf_net382));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net382 (.A(clknet_0_net382),
    .X(clknet_1_1__leaf_net382));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net376 (.A(net376),
    .X(clknet_0_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net376 (.A(clknet_0_net376),
    .X(clknet_1_0__leaf_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net376 (.A(clknet_0_net376),
    .X(clknet_1_1__leaf_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net129 (.A(net129),
    .X(clknet_0_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net129 (.A(clknet_0_net129),
    .X(clknet_1_0__leaf_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net129 (.A(clknet_0_net129),
    .X(clknet_1_1__leaf_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net139 (.A(net139),
    .X(clknet_0_net139));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net139 (.A(clknet_0_net139),
    .X(clknet_1_0__leaf_net139));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net139 (.A(clknet_0_net139),
    .X(clknet_1_1__leaf_net139));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net120 (.A(net120),
    .X(clknet_0_net120));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net120 (.A(clknet_0_net120),
    .X(clknet_1_0__leaf_net120));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net120 (.A(net941),
    .X(clknet_1_1__leaf_net120));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net463 (.A(net463),
    .X(clknet_0_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net463 (.A(clknet_0_net463),
    .X(clknet_1_0__leaf_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net463 (.A(clknet_0_net463),
    .X(clknet_1_1__leaf_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net515 (.A(net515),
    .X(clknet_0_net515));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net515 (.A(clknet_0_net515),
    .X(clknet_1_0__leaf_net515));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net515 (.A(clknet_0_net515),
    .X(clknet_1_1__leaf_net515));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net122 (.A(net122),
    .X(clknet_0_net122));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net122 (.A(clknet_0_net122),
    .X(clknet_1_0__leaf_net122));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net122 (.A(clknet_0_net122),
    .X(clknet_1_1__leaf_net122));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net597 (.A(net597),
    .X(clknet_0_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net597 (.A(clknet_0_net597),
    .X(clknet_1_0__leaf_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net597 (.A(clknet_0_net597),
    .X(clknet_1_1__leaf_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net127 (.A(net127),
    .X(clknet_0_net127));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net127 (.A(clknet_0_net127),
    .X(clknet_1_0__leaf_net127));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net127 (.A(clknet_0_net127),
    .X(clknet_1_1__leaf_net127));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net125 (.A(net125),
    .X(clknet_0_net125));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net125 (.A(clknet_0_net125),
    .X(clknet_1_0__leaf_net125));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net125 (.A(clknet_0_net125),
    .X(clknet_1_1__leaf_net125));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net116 (.A(net116),
    .X(clknet_0_net116));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net116 (.A(clknet_0_net116),
    .X(clknet_1_0__leaf_net116));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net116 (.A(clknet_0_net116),
    .X(clknet_1_1__leaf_net116));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net468 (.A(net468),
    .X(clknet_0_net468));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net468 (.A(clknet_0_net468),
    .X(clknet_1_0__leaf_net468));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net468 (.A(clknet_0_net468),
    .X(clknet_1_1__leaf_net468));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net465 (.A(net465),
    .X(clknet_0_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net465 (.A(clknet_0_net465),
    .X(clknet_1_0__leaf_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net465 (.A(clknet_0_net465),
    .X(clknet_1_1__leaf_net465));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net619 (.A(net619),
    .X(clknet_0_net619));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net619 (.A(clknet_0_net619),
    .X(clknet_1_0__leaf_net619));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net619 (.A(clknet_0_net619),
    .X(clknet_1_1__leaf_net619));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net572 (.A(net572),
    .X(clknet_0_net572));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net572 (.A(clknet_0_net572),
    .X(clknet_1_0__leaf_net572));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net572 (.A(clknet_0_net572),
    .X(clknet_1_1__leaf_net572));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net112 (.A(net112),
    .X(clknet_0_net112));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net112 (.A(clknet_0_net112),
    .X(clknet_1_0__leaf_net112));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net112 (.A(clknet_0_net112),
    .X(clknet_1_1__leaf_net112));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net114 (.A(net114),
    .X(clknet_0_net114));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net114 (.A(clknet_0_net114),
    .X(clknet_1_0__leaf_net114));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net114 (.A(clknet_0_net114),
    .X(clknet_1_1__leaf_net114));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net107 (.A(net107),
    .X(clknet_0_net107));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net107 (.A(clknet_0_net107),
    .X(clknet_1_0__leaf_net107));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net107 (.A(clknet_0_net107),
    .X(clknet_1_1__leaf_net107));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net113 (.A(net113),
    .X(clknet_0_net113));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net113 (.A(clknet_0_net113),
    .X(clknet_1_0__leaf_net113));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net113 (.A(clknet_0_net113),
    .X(clknet_1_1__leaf_net113));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net239 (.A(net239),
    .X(clknet_0_net239));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net239 (.A(clknet_0_net239),
    .X(clknet_1_0__leaf_net239));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net239 (.A(clknet_0_net239),
    .X(clknet_1_1__leaf_net239));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net592 (.A(net592),
    .X(clknet_0_net592));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net592 (.A(clknet_0_net592),
    .X(clknet_1_0__leaf_net592));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net592 (.A(clknet_0_net592),
    .X(clknet_1_1__leaf_net592));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net457 (.A(net457),
    .X(clknet_0_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net457 (.A(clknet_0_net457),
    .X(clknet_1_0__leaf_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net457 (.A(clknet_0_net457),
    .X(clknet_1_1__leaf_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net119 (.A(net119),
    .X(clknet_0_net119));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net119 (.A(clknet_0_net119),
    .X(clknet_1_0__leaf_net119));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net119 (.A(clknet_0_net119),
    .X(clknet_1_1__leaf_net119));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net126 (.A(net126),
    .X(clknet_0_net126));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net126 (.A(clknet_0_net126),
    .X(clknet_1_0__leaf_net126));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net126 (.A(clknet_0_net126),
    .X(clknet_1_1__leaf_net126));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net884 (.A(net884),
    .X(clknet_0_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net884 (.A(clknet_0_net884),
    .X(clknet_1_0__leaf_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net884 (.A(clknet_0_net884),
    .X(clknet_1_1__leaf_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net170 (.A(net170),
    .X(clknet_0_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net170 (.A(clknet_0_net170),
    .X(clknet_1_0__leaf_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net170 (.A(clknet_0_net170),
    .X(clknet_1_1__leaf_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net136 (.A(net136),
    .X(clknet_0_net136));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net136 (.A(clknet_0_net136),
    .X(clknet_1_0__leaf_net136));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net136 (.A(clknet_0_net136),
    .X(clknet_1_1__leaf_net136));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net103 (.A(net103),
    .X(clknet_0_net103));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net103 (.A(net938),
    .X(clknet_1_0__leaf_net103));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net103 (.A(clknet_0_net103),
    .X(clknet_1_1__leaf_net103));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net550 (.A(net550),
    .X(clknet_0_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net550 (.A(clknet_0_net550),
    .X(clknet_1_0__leaf_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net550 (.A(clknet_0_net550),
    .X(clknet_1_1__leaf_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net560 (.A(net560),
    .X(clknet_0_net560));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net560 (.A(clknet_0_net560),
    .X(clknet_1_0__leaf_net560));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net560 (.A(clknet_0_net560),
    .X(clknet_1_1__leaf_net560));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net551 (.A(net551),
    .X(clknet_0_net551));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net551 (.A(clknet_0_net551),
    .X(clknet_1_0__leaf_net551));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net551 (.A(clknet_0_net551),
    .X(clknet_1_1__leaf_net551));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net350 (.A(net350),
    .X(clknet_0_net350));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net350 (.A(clknet_0_net350),
    .X(clknet_1_0__leaf_net350));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net350 (.A(clknet_0_net350),
    .X(clknet_1_1__leaf_net350));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net354 (.A(net354),
    .X(clknet_0_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net354 (.A(clknet_0_net354),
    .X(clknet_1_0__leaf_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net354 (.A(clknet_0_net354),
    .X(clknet_1_1__leaf_net354));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net78),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net80),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net65),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net75),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net934),
    .X(net935));
 sky130_fd_sc_hd__buf_6 rebuffer6 (.A(net902),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net936),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(clknet_0_net103),
    .X(net938));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer9 (.A(net95),
    .X(net939));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer10 (.A(net65),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(clknet_0_net120),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net905),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net942),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net942),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net912),
    .X(net945));
 sky130_fd_sc_hd__clkbuf_1 clone16 (.A(in4),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net82),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net950),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net948),
    .X(net949));
 sky130_fd_sc_hd__clkbuf_1 clone20 (.A(clk),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net914),
    .X(net951));
 sky130_fd_sc_hd__clkbuf_1 clone22 (.A(clknet_0_net268),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(clknet_0_net268),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net77),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net954),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net955),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(clknet_0_net263),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(clknet_0_net137),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(clknet_1_0__leaf_net134),
    .X(net959));
 sky130_fd_sc_hd__dlymetal6s4s_1 hold31 (.A(net85),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net540),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net461),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net990),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net736),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net47),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net338),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net783),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net668),
    .X(net969));
 sky130_fd_sc_hd__clkbuf_4 hold40 (.A(net801),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net378),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net319),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net703),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net869),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net255),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net131),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net320),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net565),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net682),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net151),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net850),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net708),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net374),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net689),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net554),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net678),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net29),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net392),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net684),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net320),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net762),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net258),
    .X(net995));
 sky130_fd_sc_hd__buf_8 max_cap1 (.A(net67),
    .X(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone20_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone16_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_X (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A1 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A2 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_X (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_SCD (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_B1_N (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_Y (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A0 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B1_N (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_X (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net103_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_X (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A0 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A0 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_X (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A4 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_X (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_RESET_B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_X (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A4 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_X (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net116_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_X (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net120_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_X (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net122_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_X (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_X (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net136_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_X (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net140_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_X (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_RESET_B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_B1_N (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_X (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A0 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_Q_N (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A3 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_Y (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold50_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_S0 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_Q (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A3 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S0 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_X (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_Y (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A3 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A3 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_X (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_X (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A3 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_SCE (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_SCE (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A3 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A4 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A3 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A0 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_SCD (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_B1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S0 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_X (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A0 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A3 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_X (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_S0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_X (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A3 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_Y (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_Y (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_S0 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_Y (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_S0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_B (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A3 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_X (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_B1_N (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_Y (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A4 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_B1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_X (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S0 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_B1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A3 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_X (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_S0 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_X (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A3 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_RESET_B (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_D (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_X (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_A3 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A3 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_X (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_SCD (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SCD (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_B (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_Y (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A3 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A0 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_B1_N (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_X (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A0 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_SCE (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A3 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A0 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_Y (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A4 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_B (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_B1_N (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_X (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_S1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A0 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S0 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_Y (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A0 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_Y (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_X (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A2 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_Y (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_S0 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A2 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A0 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A4 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_Y (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_X (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B1_N (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_X (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A3 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_SCD (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_SCE (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_X (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A3 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A0 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S0 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_S0 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_X (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_S1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_DE (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_SCE (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_X (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_D (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_X (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_X (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net239_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_X (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_S1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_Y (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_S1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A3 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net251_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_X (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net269_A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_X (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A3 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_SET_B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_X (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A0 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S0 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_X (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A0 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S0 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S0 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_SCE (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A3 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_X (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net282_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_X (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_Q (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_Q (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_Q (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_DE (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_X (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_Y (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_S0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_B1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_X (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A0 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A3 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A3 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_X (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A0 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_SET_B (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_B1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_Y (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_S1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_D (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_RESET_B (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_Y (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A0 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_SCE (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_B1_N (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_Y (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_X (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A3 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_D (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A4 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_SCD (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A3 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_SCD (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_SCE (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_X (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A0 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_SET_B (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A3 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_X (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A0 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_Y (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_Q (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_X (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A0 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A4 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_X (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A3 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A2 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_Q_N (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_B (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_Q (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_Q (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_SCD (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_SCD (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_Y (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A2 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A2 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_SCD (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A0 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_X (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A0 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_Q (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_RESET_B (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_X (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A0 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_RESET_B (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A2 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_X (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A4 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_X (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_s838_D (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_X (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_S1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A3 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A2 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A3 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_X (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_Q (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_Q (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A4 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A4 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_Y (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A0 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A2 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A3 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_X (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A2 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A2 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_B1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_B (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_X (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A4 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A3 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_Y (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_B (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A2 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_B (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_X (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_B1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A2 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_Y (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A3 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_Y (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B1 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A1 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_Y (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A2 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_B (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_Y (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_S0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_S0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_B1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_S0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_Q_N (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_S0 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_D (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A3 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A3 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_B1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A3 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A2 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_X (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A3 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A0 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S0 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_Y (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net468_A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_X (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A2 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_RESET_B (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A2 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_Y (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A3 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A1 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A2 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A2 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_SCD (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_B1_N (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_X (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A2 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_X (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A2 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_SCE (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A2 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_X (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A0 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_X (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_SCE (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_SET_B (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A2 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_X (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_A (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A1 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_SCD (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_X (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A0 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A3 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_Q (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net577_A (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_X (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_X (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_D (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_B1_N (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S0 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_Y (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire145_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_Y (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_D (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_X (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_Q (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_SCE (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_B (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_B1_N (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap137_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A3 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A0 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_Y (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_Q (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_B1_N (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_B (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_B1_N (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_B1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A4 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_Q (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold43_A (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_Q (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_B1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_S0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_X (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_s831_Q (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_B1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_B1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_s832_Q (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_SET_B (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A4 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_B1 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_SET_B (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_B1 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_s840_Q (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S0 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S0 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S1 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S1 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_s841_Q (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_s842_Q (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_s843_Q (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S0 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A3 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A3 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_DE (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_X (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A3 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_Y (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A3 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A3 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A3 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_B1_N (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A4 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_Y (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold31_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_Y (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A3 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_X (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A3 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_S0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A3 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_X (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A3 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_Y (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_Y (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_Y (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_X (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_D (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A3 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_Y (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_SCE (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_SCD (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SET_B (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_SCD (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A3 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_X (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_X (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_B (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A3 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_B1_N (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_S0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_A3 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A3 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A3 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A2 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_B1_N (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_SET_B (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A3 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S0 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A0 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A3 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_B (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_B (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_D (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_B1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A2 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A2 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B1_N (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A2 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A2 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A3 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_A4 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B1_N (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_A0 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A2 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S0 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_B1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A4 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A2 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S0 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A0 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A2 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_SCD (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S0 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A3 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_B1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A3 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A2 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_B1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_S1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_A (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A2 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_A2 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A3 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A0 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_D (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A2 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_B (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A3 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A0 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A2 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S0 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A3 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_RESET_B (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_B1_N (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_B1_N (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B1_N (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A4 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A3 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A0 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_A3 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold40_A (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A0 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A0 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A3 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_A3 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_B1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A3 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_RESET_B (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A0 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_B1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_B (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_A (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B1_N (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A2 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A2 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A0 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_D (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A0 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A2 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B1_N (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_D (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_A0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A3 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A2 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_B (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A4 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_B (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S0 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A3 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A2 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A3 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_X (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_A3 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A2 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A3 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A2 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A2 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S0 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A0 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_B (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S0 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A0 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S0 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A3 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A4 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B1_N (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S0 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A3 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A2 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A0 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A2 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_S1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A2 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A2 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S0 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_B1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_B1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A2 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A2 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A2 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B1_N (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_A3 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_B (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_B1_N (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B1_N (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_A (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_A2 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A3 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A3 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_S0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A3 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_B1_N (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_B (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A2 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A3 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_B1_N (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_B (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_B1_N (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A2 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A2 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A2 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A4 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A2 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A3 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_B1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_B1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_B (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A4 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A4 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_B1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_B (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A2 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_S0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_X (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_S1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_B1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_B1_N (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_B1_N (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_X (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_RESET_B (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_RESET_B (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A2 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A3 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_B (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A4 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_D (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A3 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_B1_N (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_X (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_SCD (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_SCE (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A2 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A2 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A3 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A3 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_B (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_X (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_A0 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A0 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A2 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A2 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_A (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_A2 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A2 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_D (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_D (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_Y (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S0 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_B (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_Y (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A3 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A2 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S0 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A4 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S0 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A3 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_Y (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S0 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A0 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A3 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A0 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_S1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A2 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A3 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_Y (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold51_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A4 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A2 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_X (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_S0 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_X (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_X (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A2 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_B1 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_SET_B (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A1 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_SCD (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_RESET_B (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A2 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_Y (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_s853_Q (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S1 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S0 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A3 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_X (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S0 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S0 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_X (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A3 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_B1_N (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_Y (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_X (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_B1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_B1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_B1_N (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A2 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_B1_N (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_X (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_X (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A1 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_X (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold44_A (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_A2 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A3 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A3 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_X (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S0 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_B1_N (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_B1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_B (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_B (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_X (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_Y (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A2 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_SCD (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A2 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_Q (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap115_A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_Y (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A3 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A2 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_RESET_B (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_X (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap143_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_SCD (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_S1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_Y (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_X (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_X (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A4 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_D (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_B1_N (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A4 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_SCE (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net890_A (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_X (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_X (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_A2 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A3 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A3 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A2 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_Y (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_X (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_S0 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A3 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S0 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_SCD (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_SET_B (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_SCD (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A3 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S0 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_D (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_RESET_B (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_X (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_S0 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_S1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_SCE (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A3 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A4 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A3 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_SCE (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_B1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap115_X (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_SCD (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A3 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A2 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_B1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_X (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S0 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_SCE (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A4 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S0 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A3 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap117_X (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_B1_N (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A2 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A0 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A3 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A3 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_X (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A2 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_SCE (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B1_N (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A3 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A3 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B1_N (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap119_X (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S0 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A3 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A0 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A3 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_S1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A4 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_X (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S0 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_B1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_B1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer12_A (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_X (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_B1_N (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_B1_N (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_X (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A3 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_RESET_B (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S0 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_B1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S0 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A2 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap125_X (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S0 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_D (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_S0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B1_N (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_B1_N (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap126_X (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A4 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_A0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_B1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_X (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A2 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_B1_N (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_B1_N (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_B1_N (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A3 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_B1_N (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_B1_N (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_B1 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A1 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_X (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A3 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_B1_N (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_A2 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S0 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_S1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_SCE (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A2 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer15_A (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_X (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_B1_N (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap134_X (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A3 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A2 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A3 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S0 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_B1 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_A3 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_X (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_SET_B (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_S1 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_D (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_S1 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_S1 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_B1 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S1 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B1 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_SET_B (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A4 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_X (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A3 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_S0 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S0 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A2 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A4 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A3 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A2 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A4 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap137_X (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_B (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_S1 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A2 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A2 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_S1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_B1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_SET_B (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_SCE (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_B1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_B1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_B1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S0 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_X (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S0 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A4 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S0 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_A1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A3 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_B1_N (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A2 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_SCE (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_X (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_B1_N (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A3 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_S0 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_B1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A4 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A4 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_B1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_SCE (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_S0 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_X (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A2 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A3 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_S0 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A2 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_B1 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A3 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A3 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_B1 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap143_X (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_S0 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A1 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap144_X (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_RESET_B (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A0 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_B1_N (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_S0 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire145_X (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A3 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A0 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_X (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A0 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A3 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_B1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_B1_N (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_S1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_X (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A3 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A4 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_SCE (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_B1_N (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_X (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A3 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_SCE (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_B (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_S1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_B1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_B1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A0 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s832_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s833_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_GATE (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s831_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_GATE (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s834_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s840_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_SLEEP_B (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s828_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s829_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s830_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s835_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s837_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s849_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s850_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s864_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s839_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s851_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s852_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s853_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s854_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s856_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s872_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s883_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s857_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s858_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s859_SLEEP_B (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s860_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s861_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s862_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s863_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s878_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s881_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s882_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A4 (.DIODE(clknet_1_0__leaf_net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_SCE (.DIODE(clknet_1_0__leaf_net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S1 (.DIODE(clknet_1_0__leaf_net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net455_X (.DIODE(clknet_1_0__leaf_net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(clknet_1_1__leaf_net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(clknet_1_1__leaf_net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(clknet_1_1__leaf_net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net455_X (.DIODE(clknet_1_1__leaf_net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S1 (.DIODE(clknet_1_1__leaf_net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(clknet_1_1__leaf_net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net863_X (.DIODE(clknet_1_1__leaf_net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_RESET_B (.DIODE(clknet_1_0__leaf_net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_D (.DIODE(clknet_1_0__leaf_net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_SCD (.DIODE(clknet_1_0__leaf_net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S0 (.DIODE(clknet_1_0__leaf_net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_D (.DIODE(clknet_1_0__leaf_net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net251_X (.DIODE(clknet_1_0__leaf_net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A2 (.DIODE(clknet_1_1__leaf_net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A2 (.DIODE(clknet_1_1__leaf_net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A3 (.DIODE(clknet_1_1__leaf_net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net230_X (.DIODE(clknet_1_1__leaf_net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A0 (.DIODE(clknet_1_0__leaf_net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A3 (.DIODE(clknet_1_0__leaf_net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_SCD (.DIODE(clknet_1_0__leaf_net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_S0 (.DIODE(clknet_1_0__leaf_net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_S0 (.DIODE(clknet_1_0__leaf_net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net233_X (.DIODE(clknet_1_0__leaf_net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_RESET_B (.DIODE(clknet_1_1__leaf_net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_A1 (.DIODE(clknet_1_1__leaf_net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net233_X (.DIODE(clknet_1_1__leaf_net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A1 (.DIODE(clknet_1_1__leaf_net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A1 (.DIODE(clknet_1_1__leaf_net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net117_X (.DIODE(clknet_1_1__leaf_net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A1 (.DIODE(clknet_1_1__leaf_net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A1 (.DIODE(clknet_1_1__leaf_net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S1 (.DIODE(clknet_1_1__leaf_net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(clknet_1_1__leaf_net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net140_X (.DIODE(clknet_1_1__leaf_net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A1 (.DIODE(clknet_1_1__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A2 (.DIODE(clknet_1_1__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A2 (.DIODE(clknet_1_1__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net142_X (.DIODE(clknet_1_1__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A1 (.DIODE(clknet_1_0__leaf_net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A2 (.DIODE(clknet_1_0__leaf_net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A3 (.DIODE(clknet_1_0__leaf_net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A3 (.DIODE(clknet_1_0__leaf_net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S1 (.DIODE(clknet_1_0__leaf_net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A1 (.DIODE(clknet_1_0__leaf_net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net268_X (.DIODE(clknet_1_0__leaf_net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A3 (.DIODE(clknet_1_1__leaf_net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S0 (.DIODE(clknet_1_1__leaf_net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S1 (.DIODE(clknet_1_1__leaf_net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A4 (.DIODE(clknet_1_1__leaf_net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(clknet_1_1__leaf_net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_B1 (.DIODE(clknet_1_1__leaf_net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(clknet_1_1__leaf_net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(clknet_1_1__leaf_net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net268_X (.DIODE(clknet_1_1__leaf_net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A1 (.DIODE(clknet_1_1__leaf_net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A1 (.DIODE(clknet_1_1__leaf_net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A1 (.DIODE(clknet_1_1__leaf_net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net129_X (.DIODE(clknet_1_1__leaf_net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A1 (.DIODE(clknet_1_0__leaf_net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A3 (.DIODE(clknet_1_0__leaf_net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A3 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S0 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net120_X (.DIODE(clknet_1_0__leaf_net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_B1 (.DIODE(clknet_1_1__leaf_net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S0 (.DIODE(clknet_1_1__leaf_net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A3 (.DIODE(clknet_1_1__leaf_net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A2 (.DIODE(clknet_1_1__leaf_net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S0 (.DIODE(clknet_1_1__leaf_net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net120_X (.DIODE(clknet_1_1__leaf_net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A1 (.DIODE(clknet_1_0__leaf_net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_B1_N (.DIODE(clknet_1_0__leaf_net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A3 (.DIODE(clknet_1_0__leaf_net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(clknet_1_0__leaf_net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_RESET_B (.DIODE(clknet_1_0__leaf_net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S1 (.DIODE(clknet_1_0__leaf_net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net122_X (.DIODE(clknet_1_0__leaf_net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(clknet_1_1__leaf_net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_SCE (.DIODE(clknet_1_1__leaf_net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(clknet_1_1__leaf_net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(clknet_1_1__leaf_net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net122_X (.DIODE(clknet_1_1__leaf_net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A3 (.DIODE(clknet_1_0__leaf_net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A2 (.DIODE(clknet_1_0__leaf_net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_B1 (.DIODE(clknet_1_0__leaf_net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_SET_B (.DIODE(clknet_1_0__leaf_net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_B1 (.DIODE(clknet_1_0__leaf_net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S0 (.DIODE(clknet_1_0__leaf_net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A2 (.DIODE(clknet_1_0__leaf_net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A0 (.DIODE(clknet_1_0__leaf_net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net465_X (.DIODE(clknet_1_0__leaf_net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A1 (.DIODE(clknet_1_0__leaf_net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A3 (.DIODE(clknet_1_0__leaf_net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A1 (.DIODE(clknet_1_0__leaf_net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net112_X (.DIODE(clknet_1_0__leaf_net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A2 (.DIODE(clknet_1_1__leaf_net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A0 (.DIODE(clknet_1_1__leaf_net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A4 (.DIODE(clknet_1_1__leaf_net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net112_X (.DIODE(clknet_1_1__leaf_net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B1 (.DIODE(clknet_1_1__leaf_net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A1 (.DIODE(clknet_1_1__leaf_net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net114_X (.DIODE(clknet_1_1__leaf_net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A3 (.DIODE(clknet_1_0__leaf_net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_B1_N (.DIODE(clknet_1_0__leaf_net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A3 (.DIODE(clknet_1_0__leaf_net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net239_X (.DIODE(clknet_1_0__leaf_net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(clknet_1_1__leaf_net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(clknet_1_1__leaf_net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net136_X (.DIODE(clknet_1_1__leaf_net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_B1_N (.DIODE(clknet_1_0__leaf_net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A4 (.DIODE(clknet_1_0__leaf_net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_B1 (.DIODE(clknet_1_0__leaf_net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A3 (.DIODE(clknet_1_0__leaf_net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S0 (.DIODE(clknet_1_0__leaf_net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_S0 (.DIODE(clknet_1_0__leaf_net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net103_X (.DIODE(clknet_1_0__leaf_net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(clknet_1_1__leaf_net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A3 (.DIODE(clknet_1_1__leaf_net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A0 (.DIODE(clknet_1_1__leaf_net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(clknet_1_1__leaf_net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S0 (.DIODE(clknet_1_1__leaf_net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A1 (.DIODE(clknet_1_1__leaf_net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net103_X (.DIODE(clknet_1_1__leaf_net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_SCE (.DIODE(clknet_1_0__leaf_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A2 (.DIODE(clknet_1_0__leaf_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A3 (.DIODE(clknet_1_0__leaf_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A2 (.DIODE(clknet_1_0__leaf_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A2 (.DIODE(clknet_1_0__leaf_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_A2 (.DIODE(clknet_1_0__leaf_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net354_X (.DIODE(clknet_1_0__leaf_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_SET_B (.DIODE(clknet_1_1__leaf_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S0 (.DIODE(clknet_1_1__leaf_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(clknet_1_1__leaf_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net354_X (.DIODE(clknet_1_1__leaf_net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_X (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_B1_N (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A3 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer6_X (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer15_X (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S0 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone16_X (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer19_A (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer18_X (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer18_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone20_X (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A4 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_SCE (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_SCE (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A3 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone22_X (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold31_X (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_SCE (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold37_X (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_SET_B (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_A (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A2 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold40_X (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_S1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold43_X (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_S0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold50_X (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S0 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold56_X (.DIODE(net986));
 sky130_fd_sc_hd__xnor2_1 clone1 (.A(net992),
    .B(net906),
    .Y(net988));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net78),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer20 (.A(net100),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net994),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(net907),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer31 (.A(net997),
    .X(net998));
 sky130_fd_sc_hd__buf_6 rebuffer32 (.A(net65),
    .X(net999));
 sky130_fd_sc_hd__clkbuf_1 clone33 (.A(in0),
    .X(net1000));
 sky130_fd_sc_hd__clkbuf_1 clone34 (.A(in0),
    .X(net1001));
 sky130_fd_sc_hd__clkbuf_1 clone35 (.A(net71),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer36 (.A(clknet_1_0__leaf_net120),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer37 (.A(clknet_1_0__leaf_net120),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net793),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net810),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net784),
    .X(net1008));
 sky130_fd_sc_hd__buf_4 hold67 (.A(net792),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net838),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net13),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(in61),
    .X(net1012));
 sky130_fd_sc_hd__buf_4 hold71 (.A(net970),
    .X(net1013));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
