module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in3,
    in4,
    in5,
    in6,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out3,
    out4,
    out5,
    out6,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in3;
 input in4;
 input in5;
 input in6;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out3;
 output out4;
 output out5;
 output out6;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_0_net759;
 wire clknet_1_0__leaf_net759;
 wire clknet_1_1__leaf_net759;
 wire clknet_0_net176;
 wire clknet_1_0__leaf_net176;
 wire clknet_1_1__leaf_net176;
 wire clknet_0_net174;
 wire clknet_1_0__leaf_net174;
 wire clknet_1_1__leaf_net174;
 wire clknet_0_net758;
 wire clknet_1_0__leaf_net758;
 wire clknet_1_1__leaf_net758;
 wire clknet_0_net400;
 wire clknet_1_0__leaf_net400;
 wire clknet_1_1__leaf_net400;
 wire clknet_0_net401;
 wire clknet_1_0__leaf_net401;
 wire clknet_1_1__leaf_net401;
 wire clknet_0_net421;
 wire clknet_1_0__leaf_net421;
 wire clknet_1_1__leaf_net421;
 wire clknet_0_net398;
 wire clknet_1_0__leaf_net398;
 wire clknet_1_1__leaf_net398;
 wire clknet_0_net269;
 wire clknet_1_0__leaf_net269;
 wire clknet_1_1__leaf_net269;
 wire clknet_0_net757;
 wire clknet_1_0__leaf_net757;
 wire clknet_1_1__leaf_net757;
 wire clknet_0_net250;
 wire clknet_1_0__leaf_net250;
 wire clknet_1_1__leaf_net250;
 wire clknet_0_net827;
 wire clknet_1_0__leaf_net827;
 wire clknet_1_1__leaf_net827;
 wire clknet_0_net205;
 wire clknet_1_0__leaf_net205;
 wire clknet_1_1__leaf_net205;
 wire clknet_0_net103;
 wire clknet_1_0__leaf_net103;
 wire clknet_1_1__leaf_net103;
 wire clknet_0_net108;
 wire clknet_1_0__leaf_net108;
 wire clknet_1_1__leaf_net108;
 wire clknet_0_net274;
 wire clknet_1_0__leaf_net274;
 wire clknet_1_1__leaf_net274;
 wire clknet_0_net293;
 wire clknet_1_0__leaf_net293;
 wire clknet_1_1__leaf_net293;
 wire clknet_0_net280;
 wire clknet_1_0__leaf_net280;
 wire clknet_1_1__leaf_net280;
 wire clknet_0_net294;
 wire clknet_1_0__leaf_net294;
 wire clknet_1_1__leaf_net294;
 wire clknet_0_net264;
 wire clknet_1_0__leaf_net264;
 wire clknet_1_1__leaf_net264;
 wire clknet_0_net303;
 wire clknet_1_0__leaf_net303;
 wire clknet_1_1__leaf_net303;
 wire clknet_0_net443;
 wire clknet_1_0__leaf_net443;
 wire clknet_1_1__leaf_net443;
 wire clknet_0_net451;
 wire clknet_1_0__leaf_net451;
 wire clknet_1_1__leaf_net451;
 wire clknet_0_net448;
 wire clknet_1_0__leaf_net448;
 wire clknet_1_1__leaf_net448;
 wire clknet_0_net435;
 wire clknet_1_0__leaf_net435;
 wire clknet_1_1__leaf_net435;
 wire clknet_0_net272;
 wire clknet_1_0__leaf_net272;
 wire clknet_1_1__leaf_net272;
 wire clknet_0_net262;
 wire clknet_1_0__leaf_net262;
 wire clknet_1_1__leaf_net262;
 wire clknet_0_net292;
 wire clknet_1_0__leaf_net292;
 wire clknet_1_1__leaf_net292;
 wire clknet_0_net267;
 wire clknet_1_0__leaf_net267;
 wire clknet_1_1__leaf_net267;
 wire clknet_0_net521;
 wire clknet_1_0__leaf_net521;
 wire clknet_1_1__leaf_net521;
 wire clknet_0_net268;
 wire clknet_1_0__leaf_net268;
 wire clknet_1_1__leaf_net268;
 wire clknet_0_net265;
 wire clknet_1_0__leaf_net265;
 wire clknet_1_1__leaf_net265;
 wire clknet_0_net287;
 wire clknet_1_0__leaf_net287;
 wire clknet_1_1__leaf_net287;
 wire clknet_0_net139;
 wire clknet_1_0__leaf_net139;
 wire clknet_1_1__leaf_net139;
 wire clknet_0_net143;
 wire clknet_1_0__leaf_net143;
 wire clknet_1_1__leaf_net143;
 wire clknet_0_net187;
 wire clknet_1_0__leaf_net187;
 wire clknet_1_1__leaf_net187;
 wire clknet_0_net204;
 wire clknet_1_0__leaf_net204;
 wire clknet_1_1__leaf_net204;
 wire clknet_0_net202;
 wire clknet_1_0__leaf_net202;
 wire clknet_1_1__leaf_net202;
 wire clknet_0_net147;
 wire clknet_1_0__leaf_net147;
 wire clknet_1_1__leaf_net147;
 wire clknet_0_net142;
 wire clknet_1_0__leaf_net142;
 wire clknet_1_1__leaf_net142;
 wire clknet_0_net535;
 wire clknet_1_0__leaf_net535;
 wire clknet_1_1__leaf_net535;
 wire clknet_0_net279;
 wire clknet_1_0__leaf_net279;
 wire clknet_1_1__leaf_net279;
 wire clknet_0_net148;
 wire clknet_1_0__leaf_net148;
 wire clknet_1_1__leaf_net148;
 wire clknet_0_net146;
 wire clknet_1_0__leaf_net146;
 wire clknet_1_1__leaf_net146;
 wire clknet_0_net134;
 wire clknet_1_0__leaf_net134;
 wire clknet_1_1__leaf_net134;
 wire clknet_0_net154;
 wire clknet_1_0__leaf_net154;
 wire clknet_1_1__leaf_net154;
 wire clknet_0_net112;
 wire clknet_1_0__leaf_net112;
 wire clknet_1_1__leaf_net112;
 wire clknet_0_net372;
 wire clknet_1_0__leaf_net372;
 wire clknet_1_1__leaf_net372;
 wire clknet_0_net819;
 wire clknet_1_0__leaf_net819;
 wire clknet_1_1__leaf_net819;
 wire clknet_0_net234;
 wire clknet_1_0__leaf_net234;
 wire clknet_1_1__leaf_net234;
 wire clknet_0_net239;
 wire clknet_1_0__leaf_net239;
 wire clknet_1_1__leaf_net239;
 wire clknet_0_net233;
 wire clknet_1_0__leaf_net233;
 wire clknet_1_1__leaf_net233;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net838;
 wire net839;
 wire net840;

 sky130_fd_sc_hd__dlrbp_1 c100 (.D(net85),
    .GATE(clknet_leaf_24_clk),
    .RESET_B(net885),
    .Q(net86));
 sky130_fd_sc_hd__sdfrbp_1 c101 (.CLK(clknet_leaf_24_clk),
    .D(net891),
    .RESET_B(net77),
    .SCD(net85),
    .SCE(net69),
    .Q(net88),
    .Q_N(net87));
 sky130_fd_sc_hd__dlrtn_1 c102 (.D(net82),
    .GATE_N(clknet_leaf_24_clk),
    .RESET_B(net901),
    .Q(net89));
 sky130_fd_sc_hd__xnor2_1 c103 (.A(net948),
    .B(net87),
    .Y(net90));
 sky130_fd_sc_hd__sdfrtn_1 c104 (.CLK_N(clknet_leaf_24_clk),
    .D(net88),
    .RESET_B(net85),
    .SCD(net948),
    .SCE(net70),
    .Q(net91));
 sky130_fd_sc_hd__a21bo_1 c105 (.A1(net790),
    .A2(net66),
    .B1_N(net834),
    .X(net92));
 sky130_fd_sc_hd__xnor2_2 c106 (.A(net24),
    .B(net70),
    .Y(net93));
 sky130_fd_sc_hd__xnor2_1 c107 (.A(net68),
    .B(net795),
    .Y(net94));
 sky130_fd_sc_hd__clkbuf_1 c108 (.A(net37),
    .X(net95));
 sky130_fd_sc_hd__xnor2_1 c109 (.A(net39),
    .B(net66),
    .Y(net96));
 sky130_fd_sc_hd__dlrtn_1 c110 (.D(net92),
    .GATE_N(clknet_leaf_24_clk),
    .RESET_B(net879),
    .Q(net97));
 sky130_fd_sc_hd__dlrtn_1 c111 (.D(net96),
    .GATE_N(clknet_leaf_24_clk),
    .RESET_B(net67),
    .Q(net98));
 sky130_fd_sc_hd__clkbuf_1 c112 (.A(net734),
    .X(net99));
 sky130_fd_sc_hd__xnor2_1 c113 (.A(net37),
    .B(net91),
    .Y(net100));
 sky130_fd_sc_hd__dlrtp_1 c114 (.D(net95),
    .GATE(clknet_leaf_24_clk),
    .RESET_B(net931),
    .Q(net101));
 sky130_fd_sc_hd__clkbuf_1 c115 (.A(net67),
    .X(net102));
 sky130_fd_sc_hd__xnor2_1 c116 (.A(net98),
    .B(clknet_1_1__leaf_net757),
    .Y(net103));
 sky130_fd_sc_hd__dlrtp_1 c117 (.D(net0),
    .GATE(clknet_leaf_21_clk),
    .RESET_B(clknet_1_1__leaf_net103),
    .Q(net814));
 sky130_fd_sc_hd__xnor2_1 c118 (.A(net31),
    .B(clknet_1_0__leaf_net103),
    .Y(net104));
 sky130_fd_sc_hd__sdfbbn_1 c119 (.CLK_N(clknet_leaf_24_clk),
    .D(net102),
    .RESET_B(net0),
    .SCD(net67),
    .SCE(net96),
    .SET_B(clknet_1_0__leaf_net103),
    .Q(net820),
    .Q_N(net105));
 sky130_fd_sc_hd__buf_6 c120 (.A(net734),
    .X(net106));
 sky130_fd_sc_hd__dlrtp_1 c121 (.D(net100),
    .GATE(clknet_leaf_22_clk),
    .RESET_B(net31),
    .Q(net107));
 sky130_fd_sc_hd__xnor2_1 c122 (.A(net104),
    .B(net93),
    .Y(net108));
 sky130_fd_sc_hd__edfxbp_1 c123 (.CLK(clknet_leaf_23_clk),
    .D(clknet_1_1__leaf_net108),
    .DE(net94),
    .Q(net110),
    .Q_N(net109));
 sky130_fd_sc_hd__edfxtp_1 c124 (.CLK(clknet_leaf_23_clk),
    .D(net99),
    .DE(clknet_1_0__leaf_net108),
    .Q(net111));
 sky130_fd_sc_hd__sdlclkp_1 c125 (.CLK(clknet_leaf_22_clk),
    .GATE(net97),
    .SCE(net95),
    .GCLK(net112));
 sky130_fd_sc_hd__buf_4 c126 (.A(in14),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_4 c127 (.A(net113),
    .X(net114));
 sky130_fd_sc_hd__buf_1 c128 (.A(net803),
    .X(net115));
 sky130_fd_sc_hd__buf_1 c129 (.A(net804),
    .X(net116));
 sky130_fd_sc_hd__xnor2_4 c130 (.A(net806),
    .B(net795),
    .Y(net117));
 sky130_fd_sc_hd__buf_2 c131 (.A(in14),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_4 c132 (.A(net117),
    .X(net119));
 sky130_fd_sc_hd__buf_4 c133 (.A(net794),
    .X(net120));
 sky130_fd_sc_hd__buf_2 c134 (.A(net116),
    .X(net121));
 sky130_fd_sc_hd__xnor2_4 c135 (.A(net806),
    .B(net120),
    .Y(net122));
 sky130_fd_sc_hd__xnor2_2 c136 (.A(net121),
    .B(net120),
    .Y(net123));
 sky130_fd_sc_hd__buf_1 c137 (.A(net115),
    .X(net124));
 sky130_fd_sc_hd__mux4_2 c138 (.A0(net116),
    .A1(net803),
    .A2(net788),
    .A3(net113),
    .S0(net119),
    .S1(net836),
    .X(net125));
 sky130_fd_sc_hd__sdfxbp_1 c139 (.CLK(clknet_leaf_33_clk),
    .D(net123),
    .SCD(net117),
    .SCE(net805),
    .Q(net127),
    .Q_N(net126));
 sky130_fd_sc_hd__buf_1 c140 (.A(net749),
    .X(net128));
 sky130_fd_sc_hd__mux4_1 c141 (.A0(net124),
    .A1(net125),
    .A2(net123),
    .A3(net836),
    .S0(net114),
    .S1(net116),
    .X(net129));
 sky130_fd_sc_hd__xnor2_1 c142 (.A(net119),
    .B(net115),
    .Y(net130));
 sky130_fd_sc_hd__clkbuf_2 c143 (.A(net748),
    .X(net131));
 sky130_fd_sc_hd__xnor2_4 c144 (.A(net797),
    .B(net120),
    .Y(net132));
 sky130_fd_sc_hd__xnor2_1 c145 (.A(net132),
    .B(net806),
    .Y(net133));
 sky130_fd_sc_hd__sdlclkp_2 c146 (.CLK(clknet_leaf_33_clk),
    .GATE(net130),
    .SCE(net133),
    .GCLK(net134));
 sky130_fd_sc_hd__clkbuf_8 c147 (.A(net751),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 c148 (.A(net750),
    .X(net136));
 sky130_fd_sc_hd__xnor2_4 c149 (.A(net803),
    .B(net756),
    .Y(net137));
 sky130_fd_sc_hd__xnor2_4 c150 (.A(net807),
    .B(net126),
    .Y(net138));
 sky130_fd_sc_hd__sdlclkp_4 c151 (.CLK(clknet_leaf_32_clk),
    .GATE(net8),
    .SCE(net122),
    .GCLK(net139));
 sky130_fd_sc_hd__xnor2_4 c152 (.A(net2),
    .B(net138),
    .Y(net140));
 sky130_fd_sc_hd__xnor2_2 c153 (.A(net800),
    .B(net137),
    .Y(net141));
 sky130_fd_sc_hd__xnor2_1 c154 (.A(net137),
    .B(clknet_1_1__leaf_net139),
    .Y(net142));
 sky130_fd_sc_hd__xnor2_1 c155 (.A(clknet_1_0__leaf_net139),
    .B(net127),
    .Y(net143));
 sky130_fd_sc_hd__xnor2_2 c156 (.A(net127),
    .B(net128),
    .Y(net144));
 sky130_fd_sc_hd__xnor2_2 c157 (.A(net138),
    .B(net144),
    .Y(net145));
 sky130_fd_sc_hd__xnor2_1 c158 (.A(net138),
    .B(clknet_1_0__leaf_net142),
    .Y(net146));
 sky130_fd_sc_hd__a21bo_1 c159 (.A1(net141),
    .A2(net138),
    .B1_N(clknet_1_0__leaf_net143),
    .X(net147));
 sky130_fd_sc_hd__xnor2_1 c160 (.A(net144),
    .B(clknet_1_0__leaf_net142),
    .Y(net148));
 sky130_fd_sc_hd__dfrbp_2 c161 (.CLK(clknet_leaf_30_clk),
    .D(clknet_1_1__leaf_net148),
    .RESET_B(clknet_1_1__leaf_net147),
    .Q(net150),
    .Q_N(net149));
 sky130_fd_sc_hd__a21bo_4 c162 (.A1(net807),
    .A2(net145),
    .B1_N(net942),
    .X(net151));
 sky130_fd_sc_hd__sdfxbp_1 c163 (.CLK(clknet_leaf_32_clk),
    .D(net128),
    .SCD(clknet_1_0__leaf_net139),
    .SCE(clknet_1_0__leaf_net147),
    .Q(net153),
    .Q_N(net152));
 sky130_fd_sc_hd__a21bo_1 c164 (.A1(net136),
    .A2(clknet_1_1__leaf_net134),
    .B1_N(net140),
    .X(net154));
 sky130_fd_sc_hd__sdfxtp_1 c165 (.CLK(clknet_leaf_32_clk),
    .D(clknet_1_0__leaf_net147),
    .SCD(net137),
    .SCE(clknet_1_0__leaf_net154),
    .Q(net155));
 sky130_fd_sc_hd__sdfxtp_1 c166 (.CLK(clknet_leaf_32_clk),
    .D(net10),
    .SCD(net8),
    .SCE(net917),
    .Q(net156));
 sky130_fd_sc_hd__sdfxtp_2 c167 (.CLK(clknet_leaf_30_clk),
    .D(net875),
    .SCD(clknet_1_1__leaf_net147),
    .SCE(net897),
    .Q(net157));
 sky130_fd_sc_hd__clkbuf_1 c168 (.A(net894),
    .X(net158));
 sky130_fd_sc_hd__dfrbp_1 c169 (.CLK(clknet_leaf_31_clk),
    .D(net928),
    .RESET_B(net12),
    .Q(net160),
    .Q_N(net159));
 sky130_fd_sc_hd__xnor2_1 c170 (.A(net155),
    .B(net40),
    .Y(net161));
 sky130_fd_sc_hd__a21bo_4 c171 (.A1(net132),
    .A2(net36),
    .B1_N(net799),
    .X(net813));
 sky130_fd_sc_hd__dfrtn_1 c172 (.CLK_N(clknet_leaf_30_clk),
    .D(clknet_1_0__leaf_net148),
    .RESET_B(net122),
    .Q(net162));
 sky130_fd_sc_hd__clkbuf_4 c173 (.A(net115),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 c174 (.A(net894),
    .X(net164));
 sky130_fd_sc_hd__xnor2_1 c175 (.A(net921),
    .B(net163),
    .Y(net165));
 sky130_fd_sc_hd__dfrtp_4 c176 (.CLK(clknet_leaf_31_clk),
    .D(net28),
    .RESET_B(net151),
    .Q(net166));
 sky130_fd_sc_hd__xnor2_1 c177 (.A(net163),
    .B(net166),
    .Y(net167));
 sky130_fd_sc_hd__dfbbn_1 c178 (.CLK_N(clknet_leaf_30_clk),
    .D(net167),
    .RESET_B(net166),
    .SET_B(net26),
    .Q(net169),
    .Q_N(net168));
 sky130_fd_sc_hd__a21bo_1 c179 (.A1(net156),
    .A2(net169),
    .B1_N(net36),
    .X(net170));
 sky130_fd_sc_hd__dfrtp_1 c180 (.CLK(clknet_leaf_31_clk),
    .D(net165),
    .RESET_B(net848),
    .Q(net171));
 sky130_fd_sc_hd__mux4_1 c181 (.A0(net40),
    .A1(net15),
    .A2(net170),
    .A3(net171),
    .S0(net167),
    .S1(net132),
    .X(net172));
 sky130_fd_sc_hd__dfrtp_1 c182 (.CLK(clknet_leaf_32_clk),
    .D(net167),
    .RESET_B(clknet_1_0__leaf_net759),
    .Q(net173));
 sky130_fd_sc_hd__a21bo_1 c183 (.A1(net171),
    .A2(net163),
    .B1_N(clknet_1_1__leaf_net759),
    .X(net174));
 sky130_fd_sc_hd__a31o_1 c184 (.A1(net145),
    .A2(net171),
    .A3(net917),
    .B1(clknet_1_0__leaf_net759),
    .X(net175));
 sky130_fd_sc_hd__xnor2_1 c185 (.A(net159),
    .B(clknet_1_1__leaf_net759),
    .Y(net176));
 sky130_fd_sc_hd__a31o_1 c186 (.A1(clknet_1_0__leaf_net176),
    .A2(net168),
    .A3(net171),
    .B1(net162),
    .X(net177));
 sky130_fd_sc_hd__dfsbp_1 c187 (.CLK(clknet_leaf_31_clk),
    .D(net177),
    .SET_B(clknet_1_0__leaf_net174),
    .Q(net179),
    .Q_N(net178));
 sky130_fd_sc_hd__dfsbp_2 c188 (.CLK(clknet_leaf_31_clk),
    .D(net175),
    .SET_B(net849),
    .Q(net181),
    .Q_N(net180));
 sky130_fd_sc_hd__dfxbp_1 c189 (.CLK(clknet_leaf_27_clk),
    .D(net9),
    .Q(net183),
    .Q_N(net182));
 sky130_fd_sc_hd__xnor2_2 c190 (.A(net141),
    .B(net135),
    .Y(net184));
 sky130_fd_sc_hd__dfstp_1 c191 (.CLK(clknet_leaf_31_clk),
    .D(net165),
    .SET_B(net60),
    .Q(net185));
 sky130_fd_sc_hd__dfxtp_1 c192 (.CLK(clknet_leaf_29_clk),
    .D(net184),
    .Q(net186));
 sky130_fd_sc_hd__buf_1 c193 (.A(clknet_1_1__leaf_net143),
    .X(net187));
 sky130_fd_sc_hd__xnor2_1 c194 (.A(net179),
    .B(net183),
    .Y(net188));
 sky130_fd_sc_hd__dfstp_1 c195 (.CLK(clknet_leaf_30_clk),
    .D(net871),
    .SET_B(net0),
    .Q(net189));
 sky130_fd_sc_hd__xnor2_1 c196 (.A(net188),
    .B(net53),
    .Y(net190));
 sky130_fd_sc_hd__xnor2_4 c197 (.A(net43),
    .B(net180),
    .Y(net191));
 sky130_fd_sc_hd__dfstp_1 c198 (.CLK(clknet_leaf_27_clk),
    .D(net60),
    .SET_B(net868),
    .Q(net192));
 sky130_fd_sc_hd__dlrbn_1 c199 (.D(net918),
    .GATE_N(clknet_leaf_27_clk),
    .RESET_B(net184),
    .Q(net193));
 sky130_fd_sc_hd__xnor2_1 c200 (.A(net59),
    .B(clknet_1_0__leaf_net187),
    .Y(net194));
 sky130_fd_sc_hd__buf_1 c201 (.A(net190),
    .X(net195));
 sky130_fd_sc_hd__dlrbn_1 c202 (.D(net195),
    .GATE_N(clknet_leaf_27_clk),
    .RESET_B(net934),
    .Q(net197),
    .Q_N(net196));
 sky130_fd_sc_hd__dlrbp_2 c203 (.D(net194),
    .GATE(clknet_leaf_27_clk),
    .RESET_B(clknet_1_0__leaf_net757),
    .Q(net199),
    .Q_N(net198));
 sky130_fd_sc_hd__dlrbp_1 c204 (.D(net880),
    .GATE(clknet_leaf_27_clk),
    .RESET_B(net195),
    .Q(net200));
 sky130_fd_sc_hd__dlrtn_1 c205 (.D(clknet_1_1__leaf_net174),
    .GATE_N(clknet_leaf_27_clk),
    .RESET_B(net190),
    .Q(net201));
 sky130_fd_sc_hd__xnor2_1 c206 (.A(net193),
    .B(clknet_1_0__leaf_net187),
    .Y(net202));
 sky130_fd_sc_hd__dlrtn_1 c207 (.D(net197),
    .GATE_N(clknet_leaf_12_clk),
    .RESET_B(clknet_1_1__leaf_net202),
    .Q(net203));
 sky130_fd_sc_hd__xnor2_1 c208 (.A(net200),
    .B(clknet_1_0__leaf_net187),
    .Y(net204));
 sky130_fd_sc_hd__mux4_1 c209 (.A0(net189),
    .A1(net196),
    .A2(net198),
    .A3(net834),
    .S0(net201),
    .S1(clknet_1_0__leaf_net757),
    .X(net205));
 sky130_fd_sc_hd__xnor2_2 c210 (.A(net798),
    .B(net192),
    .Y(net206));
 sky130_fd_sc_hd__buf_1 c211 (.A(net733),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_1 c212 (.A(net732),
    .X(net208));
 sky130_fd_sc_hd__xnor2_1 c213 (.A(net79),
    .B(net70),
    .Y(net209));
 sky130_fd_sc_hd__dlrtn_1 c214 (.D(net53),
    .GATE_N(clknet_leaf_28_clk),
    .RESET_B(clknet_1_0__leaf_net204),
    .Q(net210));
 sky130_fd_sc_hd__xnor2_2 c215 (.A(net797),
    .B(net868),
    .Y(net211));
 sky130_fd_sc_hd__a21bo_1 c216 (.A1(net90),
    .A2(net834),
    .B1_N(clknet_1_1__leaf_net757),
    .X(net212));
 sky130_fd_sc_hd__dlrtp_2 c217 (.D(net206),
    .GATE(clknet_leaf_19_clk),
    .RESET_B(net151),
    .Q(net823));
 sky130_fd_sc_hd__dfbbn_1 c218 (.CLK_N(clknet_leaf_19_clk),
    .D(net212),
    .RESET_B(clknet_1_0__leaf_net202),
    .SET_B(net823),
    .Q(net214),
    .Q_N(net213));
 sky130_fd_sc_hd__xnor2_4 c219 (.A(net211),
    .B(net28),
    .Y(net215));
 sky130_fd_sc_hd__xnor2_1 c220 (.A(net210),
    .B(net835),
    .Y(net216));
 sky130_fd_sc_hd__dlrtp_2 c221 (.D(clknet_1_0__leaf_net204),
    .GATE(clknet_leaf_28_clk),
    .RESET_B(net883),
    .Q(net217));
 sky130_fd_sc_hd__dlrtp_1 c222 (.D(net208),
    .GATE(clknet_leaf_24_clk),
    .RESET_B(net215),
    .Q(net218));
 sky130_fd_sc_hd__a21bo_1 c223 (.A1(net81),
    .A2(net91),
    .B1_N(net216),
    .X(net219));
 sky130_fd_sc_hd__dfbbp_1 c224 (.CLK(clknet_leaf_27_clk),
    .D(net910),
    .RESET_B(net140),
    .SET_B(clknet_1_0__leaf_net202),
    .Q(net221),
    .Q_N(net220));
 sky130_fd_sc_hd__sdfxbp_1 c225 (.CLK(clknet_leaf_27_clk),
    .D(net216),
    .SCD(net919),
    .SCE(net215),
    .Q(net223),
    .Q_N(net222));
 sky130_fd_sc_hd__sdfxbp_1 c226 (.CLK(clknet_leaf_28_clk),
    .D(net221),
    .SCD(net949),
    .SCE(net215),
    .Q(net224));
 sky130_fd_sc_hd__xnor2_1 c227 (.A(net209),
    .B(net217),
    .Y(net225));
 sky130_fd_sc_hd__sdfbbn_2 c228 (.CLK_N(clknet_leaf_27_clk),
    .D(net192),
    .RESET_B(net119),
    .SCD(net73),
    .SCE(net222),
    .SET_B(clknet_1_1__leaf_net204),
    .Q(net227),
    .Q_N(net226));
 sky130_fd_sc_hd__xnor2_4 c229 (.A(net223),
    .B(net226),
    .Y(net228));
 sky130_fd_sc_hd__a21bo_1 c230 (.A1(net224),
    .A2(net218),
    .B1_N(net223),
    .X(net229));
 sky130_fd_sc_hd__xnor2_1 c231 (.A(net227),
    .B(net110),
    .Y(net230));
 sky130_fd_sc_hd__sdfxtp_1 c232 (.CLK(clknet_leaf_22_clk),
    .D(net70),
    .SCD(net225),
    .SCE(clknet_1_0__leaf_net112),
    .Q(net231));
 sky130_fd_sc_hd__sdfxtp_1 c233 (.CLK(clknet_leaf_22_clk),
    .D(net225),
    .SCD(net900),
    .SCE(net945),
    .Q(net232));
 sky130_fd_sc_hd__a21bo_1 c234 (.A1(net230),
    .A2(net823),
    .B1_N(clknet_1_1__leaf_net112),
    .X(net233));
 sky130_fd_sc_hd__a21bo_1 c235 (.A1(net101),
    .A2(net183),
    .B1_N(clknet_1_0__leaf_net112),
    .X(net234));
 sky130_fd_sc_hd__edfxbp_1 c236 (.CLK(clknet_leaf_23_clk),
    .D(net900),
    .DE(net215),
    .Q(net235));
 sky130_fd_sc_hd__a21bo_4 c237 (.A1(net106),
    .A2(net183),
    .B1_N(net198),
    .X(net809));
 sky130_fd_sc_hd__a21bo_1 c238 (.A1(net111),
    .A2(net183),
    .B1_N(net795),
    .X(net236));
 sky130_fd_sc_hd__a21bo_1 c239 (.A1(clknet_1_1__leaf_net234),
    .A2(clknet_1_0__leaf_net112),
    .B1_N(net217),
    .X(net819));
 sky130_fd_sc_hd__a21bo_4 c240 (.A1(net91),
    .A2(net84),
    .B1_N(net809),
    .X(net237));
 sky130_fd_sc_hd__sdfxtp_1 c241 (.CLK(clknet_leaf_22_clk),
    .D(net872),
    .SCD(net215),
    .SCE(net237),
    .Q(net238));
 sky130_fd_sc_hd__a21bo_1 c242 (.A1(net237),
    .A2(net238),
    .B1_N(clknet_1_1__leaf_net234),
    .X(net239));
 sky130_fd_sc_hd__dfbbn_1 c243 (.CLK_N(clknet_leaf_21_clk),
    .D(net231),
    .RESET_B(clknet_1_1__leaf_net239),
    .SET_B(clknet_1_1__leaf_net757),
    .Q(net241),
    .Q_N(net240));
 sky130_fd_sc_hd__dfbbn_1 c244 (.CLK_N(clknet_leaf_23_clk),
    .D(clknet_1_0__leaf_net239),
    .RESET_B(net109),
    .SET_B(clknet_1_0__leaf_net234),
    .Q(net243),
    .Q_N(net242));
 sky130_fd_sc_hd__a21bo_1 c245 (.A1(net106),
    .A2(net227),
    .B1_N(net91),
    .X(net244));
 sky130_fd_sc_hd__sdfbbp_1 c246 (.CLK(clknet_leaf_22_clk),
    .D(net135),
    .RESET_B(net70),
    .SCD(clknet_1_0__leaf_net819),
    .SCE(net963),
    .SET_B(net0),
    .Q(net246),
    .Q_N(net245));
 sky130_fd_sc_hd__mux4_1 c247 (.A0(net244),
    .A1(net246),
    .A2(net182),
    .A3(net0),
    .S0(net237),
    .S1(clknet_1_0__leaf_net234),
    .X(net247));
 sky130_fd_sc_hd__a21bo_1 c248 (.A1(net93),
    .A2(net237),
    .B1_N(net761),
    .X(net830));
 sky130_fd_sc_hd__dfbbp_1 c249 (.CLK(clknet_leaf_21_clk),
    .D(net832),
    .RESET_B(clknet_1_0__leaf_net239),
    .SET_B(net761),
    .Q(net812),
    .Q_N(net248));
 sky130_fd_sc_hd__xnor2_4 c25 (.A(net800),
    .B(net6),
    .Y(net0));
 sky130_fd_sc_hd__a21bo_1 c250 (.A1(net232),
    .A2(net101),
    .B1_N(net242),
    .X(net249));
 sky130_fd_sc_hd__a41o_1 c251 (.A1(net249),
    .A2(net245),
    .A3(net823),
    .A4(clknet_1_1__leaf_net757),
    .B1(net760),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_8 c252 (.A(net120),
    .X(net251));
 sky130_fd_sc_hd__xnor2_4 c253 (.A(net131),
    .B(net251),
    .Y(net252));
 sky130_fd_sc_hd__xnor2_4 c254 (.A(net792),
    .B(net114),
    .Y(net253));
 sky130_fd_sc_hd__xnor2_1 c255 (.A(net120),
    .B(net251),
    .Y(net254));
 sky130_fd_sc_hd__buf_4 c256 (.A(net808),
    .X(net255));
 sky130_fd_sc_hd__xnor2_2 c257 (.A(net786),
    .B(net251),
    .Y(net256));
 sky130_fd_sc_hd__clkbuf_8 c258 (.A(net735),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_4 c259 (.A(net131),
    .X(net258));
 sky130_fd_sc_hd__mux4_1 c26 (.A0(net799),
    .A1(net789),
    .A2(net800),
    .A3(net0),
    .S0(net8),
    .S1(net12),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 c260 (.A(net257),
    .X(net259));
 sky130_fd_sc_hd__buf_1 c261 (.A(net735),
    .X(net260));
 sky130_fd_sc_hd__edfxtp_1 c262 (.CLK(clknet_leaf_4_clk),
    .D(net260),
    .DE(net256),
    .Q(net261));
 sky130_fd_sc_hd__sdlclkp_1 c263 (.CLK(clknet_leaf_33_clk),
    .GATE(net259),
    .SCE(net130),
    .GCLK(net262));
 sky130_fd_sc_hd__xnor2_4 c264 (.A(net258),
    .B(net257),
    .Y(net263));
 sky130_fd_sc_hd__sdlclkp_2 c265 (.CLK(clknet_leaf_34_clk),
    .GATE(net263),
    .SCE(net254),
    .GCLK(net264));
 sky130_fd_sc_hd__xnor2_1 c266 (.A(net792),
    .B(clknet_1_0__leaf_net262),
    .Y(net265));
 sky130_fd_sc_hd__buf_2 c267 (.A(net261),
    .X(net266));
 sky130_fd_sc_hd__xnor2_1 c268 (.A(clknet_1_0__leaf_net262),
    .B(net802),
    .Y(net267));
 sky130_fd_sc_hd__xnor2_1 c269 (.A(clknet_1_0__leaf_net267),
    .B(net257),
    .Y(net268));
 sky130_fd_sc_hd__xnor2_4 c27 (.A(net801),
    .B(net17),
    .Y(net2));
 sky130_fd_sc_hd__xnor2_1 c270 (.A(clknet_1_0__leaf_net268),
    .B(clknet_1_0__leaf_net758),
    .Y(net269));
 sky130_fd_sc_hd__sdfxbp_1 c271 (.CLK(clknet_leaf_34_clk),
    .D(net133),
    .SCD(net258),
    .SCE(clknet_1_0__leaf_net268),
    .Q(net271),
    .Q_N(net270));
 sky130_fd_sc_hd__a21bo_1 c272 (.A1(clknet_1_0__leaf_net264),
    .A2(clknet_1_1__leaf_net268),
    .B1_N(clknet_1_0__leaf_net265),
    .X(net272));
 sky130_fd_sc_hd__xnor2_4 c273 (.A(net808),
    .B(net837),
    .Y(net273));
 sky130_fd_sc_hd__sdlclkp_4 c274 (.CLK(clknet_leaf_35_clk),
    .GATE(net259),
    .SCE(clknet_1_0__leaf_net272),
    .GCLK(net274));
 sky130_fd_sc_hd__dfrbp_2 c275 (.CLK(clknet_leaf_35_clk),
    .D(clknet_1_0__leaf_net146),
    .RESET_B(net787),
    .Q(net276),
    .Q_N(net275));
 sky130_fd_sc_hd__dfrbp_1 c276 (.CLK(clknet_leaf_35_clk),
    .D(net254),
    .RESET_B(net14),
    .Q(net278),
    .Q_N(net277));
 sky130_fd_sc_hd__xnor2_1 c277 (.A(net260),
    .B(clknet_1_1__leaf_net142),
    .Y(net279));
 sky130_fd_sc_hd__xnor2_1 c278 (.A(clknet_1_0__leaf_net274),
    .B(net15),
    .Y(net280));
 sky130_fd_sc_hd__dfrtn_1 c279 (.CLK_N(clknet_leaf_35_clk),
    .D(net278),
    .RESET_B(clknet_1_1__leaf_net146),
    .Q(net281));
 sky130_fd_sc_hd__buf_1 c28 (.A(net793),
    .X(net3));
 sky130_fd_sc_hd__dfrtp_4 c280 (.CLK(clknet_leaf_30_clk),
    .D(net14),
    .RESET_B(clknet_1_1__leaf_net280),
    .Q(net282));
 sky130_fd_sc_hd__dfrtp_1 c281 (.CLK(clknet_leaf_34_clk),
    .D(clknet_1_1__leaf_net272),
    .RESET_B(net842),
    .Q(net283));
 sky130_fd_sc_hd__xnor2_1 c282 (.A(net17),
    .B(net3),
    .Y(net284));
 sky130_fd_sc_hd__a21bo_1 c283 (.A1(net276),
    .A2(net284),
    .B1_N(net283),
    .X(net285));
 sky130_fd_sc_hd__dfrtp_4 c284 (.CLK(clknet_leaf_34_clk),
    .D(net256),
    .RESET_B(net273),
    .Q(net286));
 sky130_fd_sc_hd__xnor2_1 c285 (.A(clknet_1_1__leaf_net265),
    .B(net276),
    .Y(net287));
 sky130_fd_sc_hd__dfsbp_1 c286 (.CLK(clknet_leaf_35_clk),
    .D(net285),
    .SET_B(clknet_1_0__leaf_net287),
    .Q(net289),
    .Q_N(net288));
 sky130_fd_sc_hd__sdfxbp_1 c287 (.CLK(clknet_leaf_35_clk),
    .D(net284),
    .SCD(net140),
    .SCE(net285),
    .Q(net291),
    .Q_N(net290));
 sky130_fd_sc_hd__xnor2_1 c288 (.A(clknet_1_1__leaf_net262),
    .B(net277),
    .Y(net292));
 sky130_fd_sc_hd__a21bo_1 c289 (.A1(net289),
    .A2(net157),
    .B1_N(clknet_1_1__leaf_net274),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_2 c29 (.A(net785),
    .X(net4));
 sky130_fd_sc_hd__a21bo_1 c290 (.A1(net281),
    .A2(clknet_1_0__leaf_net280),
    .B1_N(clknet_1_0__leaf_net292),
    .X(net294));
 sky130_fd_sc_hd__sdfbbn_2 c291 (.CLK_N(clknet_leaf_0_clk),
    .D(net3),
    .RESET_B(clknet_1_0__leaf_net294),
    .SCD(net940),
    .SCE(clknet_1_0__leaf_net280),
    .SET_B(net277),
    .Q(net296),
    .Q_N(net295));
 sky130_fd_sc_hd__sdfbbn_2 c292 (.CLK_N(clknet_leaf_35_clk),
    .D(clknet_1_1__leaf_net292),
    .RESET_B(clknet_1_0__leaf_net280),
    .SCD(clknet_1_0__leaf_net293),
    .SCE(net285),
    .SET_B(net842),
    .Q(net298),
    .Q_N(net297));
 sky130_fd_sc_hd__sdfbbp_1 c293 (.CLK(clknet_leaf_0_clk),
    .D(net904),
    .RESET_B(clknet_1_0__leaf_net294),
    .SCD(net297),
    .SCE(net281),
    .SET_B(net756),
    .Q(net300),
    .Q_N(net299));
 sky130_fd_sc_hd__dfsbp_1 c294 (.CLK(clknet_leaf_0_clk),
    .D(net12),
    .SET_B(net2),
    .Q(net302),
    .Q_N(net301));
 sky130_fd_sc_hd__xnor2_1 c295 (.A(clknet_1_1__leaf_net264),
    .B(net301),
    .Y(net303));
 sky130_fd_sc_hd__sdfxtp_1 c296 (.CLK(clknet_leaf_30_clk),
    .D(net805),
    .SCD(net29),
    .SCE(net813),
    .Q(net304));
 sky130_fd_sc_hd__a31o_1 c297 (.A1(net170),
    .A2(net886),
    .A3(net799),
    .B1(net848),
    .X(net305));
 sky130_fd_sc_hd__sdfxtp_1 c298 (.CLK(clknet_leaf_0_clk),
    .D(net305),
    .SCD(net286),
    .SCE(net163),
    .Q(net306));
 sky130_fd_sc_hd__a21bo_2 c299 (.A1(net169),
    .A2(net856),
    .B1_N(net34),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_2 c30 (.A(net4),
    .X(net5));
 sky130_fd_sc_hd__a21bo_1 c300 (.A1(net164),
    .A2(net140),
    .B1_N(net298),
    .X(net308));
 sky130_fd_sc_hd__dfstp_1 c301 (.CLK(clknet_leaf_30_clk),
    .D(net158),
    .SET_B(net308),
    .Q(net309));
 sky130_fd_sc_hd__xnor2_1 c302 (.A(clknet_1_1__leaf_net280),
    .B(net168),
    .Y(net310));
 sky130_fd_sc_hd__dfstp_2 c303 (.CLK(clknet_leaf_1_clk),
    .D(net308),
    .SET_B(net163),
    .Q(net311));
 sky130_fd_sc_hd__dfstp_2 c304 (.CLK(clknet_leaf_0_clk),
    .D(clknet_1_1__leaf_net268),
    .SET_B(net887),
    .Q(net312));
 sky130_fd_sc_hd__dlrbn_1 c305 (.D(net933),
    .GATE_N(clknet_leaf_12_clk),
    .RESET_B(net308),
    .Q(net314),
    .Q_N(net313));
 sky130_fd_sc_hd__xnor2_2 c306 (.A(net15),
    .B(net311),
    .Y(net315));
 sky130_fd_sc_hd__dlrbn_1 c307 (.D(net922),
    .GATE_N(clknet_leaf_0_clk),
    .RESET_B(net151),
    .Q(net316));
 sky130_fd_sc_hd__mux4_1 c308 (.A0(net959),
    .A1(net282),
    .A2(net161),
    .A3(net273),
    .S0(net312),
    .S1(net36),
    .X(net317));
 sky130_fd_sc_hd__xnor2_4 c309 (.A(net315),
    .B(net149),
    .Y(net318));
 sky130_fd_sc_hd__clkbuf_4 c31 (.A(net3),
    .X(net6));
 sky130_fd_sc_hd__dlrbp_1 c310 (.D(net309),
    .GATE(clknet_leaf_29_clk),
    .RESET_B(net308),
    .Q(net319));
 sky130_fd_sc_hd__sdfbbn_1 c311 (.CLK_N(clknet_leaf_29_clk),
    .D(net317),
    .RESET_B(net312),
    .SCD(net308),
    .SCE(net166),
    .SET_B(net304),
    .Q(net321),
    .Q_N(net320));
 sky130_fd_sc_hd__xnor2_2 c312 (.A(net319),
    .B(net311),
    .Y(net322));
 sky130_fd_sc_hd__a21bo_1 c313 (.A1(net161),
    .A2(net322),
    .B1_N(net321),
    .X(net323));
 sky130_fd_sc_hd__dlrbp_1 c314 (.D(net323),
    .GATE(clknet_leaf_29_clk),
    .RESET_B(net318),
    .Q(net324));
 sky130_fd_sc_hd__dlrtn_1 c315 (.D(net286),
    .GATE_N(clknet_leaf_18_clk),
    .RESET_B(net51),
    .Q(net325));
 sky130_fd_sc_hd__dlrtn_1 c316 (.D(net252),
    .GATE_N(clknet_leaf_29_clk),
    .RESET_B(net122),
    .Q(net326));
 sky130_fd_sc_hd__xnor2_1 c317 (.A(net201),
    .B(net312),
    .Y(net327));
 sky130_fd_sc_hd__xnor2_1 c318 (.A(net788),
    .B(net27),
    .Y(net328));
 sky130_fd_sc_hd__sdfxtp_1 c319 (.CLK(clknet_leaf_29_clk),
    .D(net843),
    .SCD(net36),
    .SCE(clknet_1_1__leaf_net294),
    .Q(net329));
 sky130_fd_sc_hd__buf_2 c32 (.A(net4),
    .X(net7));
 sky130_fd_sc_hd__dlrtn_1 c320 (.D(net184),
    .GATE_N(clknet_leaf_29_clk),
    .RESET_B(net296),
    .Q(net330));
 sky130_fd_sc_hd__dlrtp_1 c321 (.D(net51),
    .GATE(clknet_leaf_29_clk),
    .RESET_B(net328),
    .Q(net331));
 sky130_fd_sc_hd__dfbbn_1 c322 (.CLK_N(clknet_leaf_29_clk),
    .D(net173),
    .RESET_B(clknet_1_0__leaf_net205),
    .SET_B(net843),
    .Q(net332));
 sky130_fd_sc_hd__dlrtp_1 c323 (.D(net865),
    .GATE(clknet_leaf_29_clk),
    .RESET_B(clknet_1_0__leaf_net205),
    .Q(net333));
 sky130_fd_sc_hd__xnor2_1 c324 (.A(net798),
    .B(net962),
    .Y(net334));
 sky130_fd_sc_hd__dlrtp_1 c325 (.D(clknet_1_1__leaf_net176),
    .GATE(clknet_leaf_30_clk),
    .RESET_B(net252),
    .Q(net335));
 sky130_fd_sc_hd__a21bo_1 c326 (.A1(net333),
    .A2(net334),
    .B1_N(net312),
    .X(net336));
 sky130_fd_sc_hd__xnor2_1 c327 (.A(net332),
    .B(net335),
    .Y(net337));
 sky130_fd_sc_hd__xnor2_4 c328 (.A(net324),
    .B(net286),
    .Y(net338));
 sky130_fd_sc_hd__xnor2_2 c329 (.A(net335),
    .B(net338),
    .Y(net339));
 sky130_fd_sc_hd__xnor2_2 c33 (.A(net6),
    .B(net10),
    .Y(net8));
 sky130_fd_sc_hd__xnor2_1 c330 (.A(net330),
    .B(net338),
    .Y(net340));
 sky130_fd_sc_hd__mux4_1 c331 (.A0(net340),
    .A1(net286),
    .A2(net27),
    .A3(net338),
    .S0(net318),
    .S1(net330),
    .X(net341));
 sky130_fd_sc_hd__dfbbn_1 c332 (.CLK_N(clknet_leaf_29_clk),
    .D(net336),
    .RESET_B(net51),
    .SET_B(net338),
    .Q(net343),
    .Q_N(net342));
 sky130_fd_sc_hd__dfbbp_1 c333 (.CLK(clknet_leaf_29_clk),
    .D(net343),
    .RESET_B(net318),
    .SET_B(net862),
    .Q(net344));
 sky130_fd_sc_hd__a21bo_1 c334 (.A1(net334),
    .A2(net342),
    .B1_N(net338),
    .X(net345));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(net329),
    .A1(net340),
    .A2(net339),
    .A3(net338),
    .S0(net26),
    .S1(clknet_1_0__leaf_net202),
    .X(net346));
 sky130_fd_sc_hd__xnor2_1 c336 (.A(net46),
    .B(net282),
    .Y(net347));
 sky130_fd_sc_hd__edfxbp_1 c337 (.CLK(clknet_leaf_25_clk),
    .D(net71),
    .DE(net74),
    .Q(net348));
 sky130_fd_sc_hd__edfxtp_1 c338 (.CLK(clknet_leaf_28_clk),
    .D(clknet_1_1__leaf_net205),
    .DE(net298),
    .Q(net349));
 sky130_fd_sc_hd__clkbuf_1 c339 (.A(net228),
    .X(net350));
 sky130_fd_sc_hd__xnor2_4 c34 (.A(net7),
    .B(net791),
    .Y(net9));
 sky130_fd_sc_hd__sdlclkp_1 c340 (.CLK(clknet_leaf_22_clk),
    .GATE(net214),
    .SCE(clknet_1_0__leaf_net202),
    .GCLK(net351));
 sky130_fd_sc_hd__sdfxbp_1 c341 (.CLK(clknet_leaf_19_clk),
    .D(net351),
    .SCD(net71),
    .SCE(net229),
    .Q(net352));
 sky130_fd_sc_hd__xnor2_1 c342 (.A(net326),
    .B(net295),
    .Y(net353));
 sky130_fd_sc_hd__dlymetal6s2s_1 c343 (.A(net953),
    .X(net354));
 sky130_fd_sc_hd__xnor2_4 c344 (.A(net786),
    .B(net228),
    .Y(net355));
 sky130_fd_sc_hd__xnor2_1 c345 (.A(net325),
    .B(net355),
    .Y(net356));
 sky130_fd_sc_hd__xnor2_1 c346 (.A(net353),
    .B(net45),
    .Y(net357));
 sky130_fd_sc_hd__sdfxbp_1 c347 (.CLK(clknet_leaf_19_clk),
    .D(net902),
    .SCD(net228),
    .SCE(clknet_1_0__leaf_net202),
    .Q(net358));
 sky130_fd_sc_hd__xnor2_1 c348 (.A(net282),
    .B(net213),
    .Y(net359));
 sky130_fd_sc_hd__xnor2_4 c349 (.A(net355),
    .B(net354),
    .Y(net360));
 sky130_fd_sc_hd__xnor2_4 c35 (.A(net791),
    .B(net794),
    .Y(net10));
 sky130_fd_sc_hd__xnor2_1 c350 (.A(net75),
    .B(net46),
    .Y(net361));
 sky130_fd_sc_hd__a21bo_2 c351 (.A1(net347),
    .A2(net295),
    .B1_N(net355),
    .X(net362));
 sky130_fd_sc_hd__sdfxtp_1 c352 (.CLK(clknet_leaf_19_clk),
    .D(net361),
    .SCD(net360),
    .SCE(net362),
    .Q(net363));
 sky130_fd_sc_hd__mux4_1 c353 (.A0(net358),
    .A1(net353),
    .A2(net363),
    .A3(net355),
    .S0(net347),
    .S1(clknet_1_0__leaf_net202),
    .X(net364));
 sky130_fd_sc_hd__sdfxtp_1 c354 (.CLK(clknet_leaf_17_clk),
    .D(net69),
    .SCD(net181),
    .SCE(net765),
    .Q(net365));
 sky130_fd_sc_hd__a21bo_1 c355 (.A1(net359),
    .A2(net355),
    .B1_N(net320),
    .X(net366));
 sky130_fd_sc_hd__sdlclkp_2 c356 (.CLK(clknet_leaf_19_clk),
    .GATE(net366),
    .SCE(net347),
    .GCLK(net367));
 sky130_fd_sc_hd__sdfxtp_1 c357 (.CLK(clknet_leaf_19_clk),
    .D(net889),
    .SCD(net11),
    .SCE(net215),
    .Q(net368));
 sky130_fd_sc_hd__a21bo_1 c358 (.A1(clknet_1_1__leaf_net250),
    .A2(net368),
    .B1_N(net135),
    .X(net369));
 sky130_fd_sc_hd__xnor2_2 c359 (.A(net199),
    .B(net820),
    .Y(net829));
 sky130_fd_sc_hd__clkbuf_4 c36 (.A(net742),
    .X(net11));
 sky130_fd_sc_hd__a21bo_1 c360 (.A1(net357),
    .A2(net199),
    .B1_N(net113),
    .X(net370));
 sky130_fd_sc_hd__a31o_1 c361 (.A1(clknet_1_1__leaf_net103),
    .A2(net368),
    .A3(net840),
    .B1(net257),
    .X(net371));
 sky130_fd_sc_hd__a41o_1 c362 (.A1(net350),
    .A2(net13),
    .A3(net105),
    .A4(clknet_1_0__leaf_net233),
    .B1(clknet_1_1__leaf_net112),
    .X(net372));
 sky130_fd_sc_hd__xnor2_2 c363 (.A(net241),
    .B(net907),
    .Y(net373));
 sky130_fd_sc_hd__a21bo_1 c364 (.A1(net243),
    .A2(net373),
    .B1_N(net907),
    .X(net374));
 sky130_fd_sc_hd__xnor2_1 c365 (.A(net838),
    .B(net84),
    .Y(net375));
 sky130_fd_sc_hd__sdlclkp_4 c366 (.CLK(clknet_leaf_21_clk),
    .GATE(net369),
    .SCE(net908),
    .GCLK(net376));
 sky130_fd_sc_hd__dfrbp_1 c367 (.CLK(clknet_leaf_19_clk),
    .D(net119),
    .RESET_B(net215),
    .Q(net377));
 sky130_fd_sc_hd__a41o_1 c368 (.A1(net321),
    .A2(net814),
    .A3(net83),
    .A4(net374),
    .B1(clknet_1_0__leaf_net250),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 c369 (.A0(net377),
    .A1(net376),
    .A2(net240),
    .A3(net373),
    .S0(net838),
    .S1(clknet_1_0__leaf_net112),
    .X(net827));
 sky130_fd_sc_hd__xnor2_4 c37 (.A(net6),
    .B(net10),
    .Y(net12));
 sky130_fd_sc_hd__a21bo_1 c370 (.A1(clknet_1_1__leaf_net112),
    .A2(net217),
    .B1_N(net373),
    .X(net379));
 sky130_fd_sc_hd__a31o_1 c371 (.A1(net371),
    .A2(net374),
    .A3(net320),
    .B1(clknet_1_1__leaf_net112),
    .X(net380));
 sky130_fd_sc_hd__a21bo_1 c372 (.A1(net296),
    .A2(net379),
    .B1_N(net832),
    .X(net833));
 sky130_fd_sc_hd__dfbbn_1 c373 (.CLK_N(clknet_leaf_21_clk),
    .D(net370),
    .RESET_B(net375),
    .SET_B(net374),
    .Q(net811));
 sky130_fd_sc_hd__a21bo_1 c374 (.A1(net84),
    .A2(net838),
    .B1_N(net368),
    .X(net381));
 sky130_fd_sc_hd__xnor2_1 c375 (.A(net374),
    .B(net373),
    .Y(net382));
 sky130_fd_sc_hd__dfrbp_1 c376 (.CLK(clknet_leaf_20_clk),
    .D(net380),
    .RESET_B(net382),
    .Q(net383));
 sky130_fd_sc_hd__dfbbn_1 c377 (.CLK_N(clknet_leaf_20_clk),
    .D(net381),
    .RESET_B(net383),
    .SET_B(clknet_1_1__leaf_net112),
    .Q(net385),
    .Q_N(net384));
 sky130_fd_sc_hd__xnor2_2 c378 (.A(net118),
    .B(net787),
    .Y(net386));
 sky130_fd_sc_hd__xnor2_4 c379 (.A(net258),
    .B(net255),
    .Y(net387));
 sky130_fd_sc_hd__clkbuf_4 c38 (.A(net742),
    .X(net13));
 sky130_fd_sc_hd__dfxtp_2 c380 (.CLK(clknet_leaf_34_clk),
    .D(clknet_1_0__leaf_net269),
    .Q(net388));
 sky130_fd_sc_hd__xnor2_1 c381 (.A(net114),
    .B(net387),
    .Y(net389));
 sky130_fd_sc_hd__xnor2_1 c382 (.A(clknet_1_0__leaf_net267),
    .B(clknet_1_0__leaf_net758),
    .Y(net390));
 sky130_fd_sc_hd__xnor2_1 c383 (.A(net251),
    .B(net263),
    .Y(net391));
 sky130_fd_sc_hd__dfrtn_1 c384 (.CLK_N(clknet_leaf_3_clk),
    .D(net391),
    .RESET_B(net255),
    .Q(net392));
 sky130_fd_sc_hd__dfbbp_1 c385 (.CLK(clknet_leaf_3_clk),
    .D(net392),
    .RESET_B(net391),
    .SET_B(net253),
    .Q(net394),
    .Q_N(net393));
 sky130_fd_sc_hd__clkbuf_2 c386 (.A(net860),
    .X(net395));
 sky130_fd_sc_hd__dfrtp_4 c387 (.CLK(clknet_leaf_4_clk),
    .D(net389),
    .RESET_B(net395),
    .Q(net396));
 sky130_fd_sc_hd__xnor2_4 c388 (.A(net396),
    .B(net270),
    .Y(net397));
 sky130_fd_sc_hd__xnor2_1 c389 (.A(net390),
    .B(net257),
    .Y(net398));
 sky130_fd_sc_hd__xnor2_1 c39 (.A(net5),
    .B(net7),
    .Y(net14));
 sky130_fd_sc_hd__dfrtp_4 c390 (.CLK(clknet_leaf_4_clk),
    .D(clknet_1_0__leaf_net398),
    .RESET_B(net114),
    .Q(net399));
 sky130_fd_sc_hd__a21bo_1 c391 (.A1(net786),
    .A2(net392),
    .B1_N(clknet_1_1__leaf_net758),
    .X(net400));
 sky130_fd_sc_hd__buf_1 c392 (.A(clknet_1_1__leaf_net400),
    .X(net401));
 sky130_fd_sc_hd__dfrtp_4 c393 (.CLK(clknet_leaf_4_clk),
    .D(net881),
    .RESET_B(clknet_1_1__leaf_net398),
    .Q(net402));
 sky130_fd_sc_hd__xnor2_1 c394 (.A(net397),
    .B(net255),
    .Y(net403));
 sky130_fd_sc_hd__xnor2_2 c395 (.A(net386),
    .B(net932),
    .Y(net404));
 sky130_fd_sc_hd__sdfxbp_2 c396 (.CLK(clknet_leaf_4_clk),
    .D(net932),
    .SCD(net121),
    .SCE(net404),
    .Q(net406),
    .Q_N(net405));
 sky130_fd_sc_hd__dfsbp_1 c397 (.CLK(clknet_leaf_34_clk),
    .D(clknet_1_0__leaf_net400),
    .SET_B(net404),
    .Q(net408),
    .Q_N(net407));
 sky130_fd_sc_hd__sdfrtp_1 c398 (.CLK(clknet_leaf_3_clk),
    .D(net403),
    .RESET_B(clknet_1_1__leaf_net401),
    .SCD(net252),
    .SCE(net387),
    .Q(net409));
 sky130_fd_sc_hd__xnor2_4 c399 (.A(net255),
    .B(net149),
    .Y(net410));
 sky130_fd_sc_hd__a21bo_4 c40 (.A1(net791),
    .A2(net785),
    .B1_N(net11),
    .X(net15));
 sky130_fd_sc_hd__xnor2_4 c400 (.A(net805),
    .B(net796),
    .Y(net411));
 sky130_fd_sc_hd__clkbuf_1 c401 (.A(net747),
    .X(net412));
 sky130_fd_sc_hd__xnor2_1 c402 (.A(net278),
    .B(net399),
    .Y(net413));
 sky130_fd_sc_hd__xnor2_4 c403 (.A(net410),
    .B(net117),
    .Y(net414));
 sky130_fd_sc_hd__xnor2_1 c404 (.A(net802),
    .B(net399),
    .Y(net415));
 sky130_fd_sc_hd__xnor2_1 c405 (.A(net399),
    .B(net395),
    .Y(net416));
 sky130_fd_sc_hd__xnor2_1 c406 (.A(net291),
    .B(net407),
    .Y(net417));
 sky130_fd_sc_hd__xnor2_1 c407 (.A(net909),
    .B(net290),
    .Y(net418));
 sky130_fd_sc_hd__a21bo_1 c408 (.A1(net417),
    .A2(net394),
    .B1_N(net411),
    .X(net419));
 sky130_fd_sc_hd__buf_1 c409 (.A(net747),
    .X(net420));
 sky130_fd_sc_hd__dfbbn_2 c41 (.CLK_N(clknet_leaf_0_clk),
    .D(net7),
    .RESET_B(net14),
    .SET_B(net13),
    .Q(net17),
    .Q_N(net16));
 sky130_fd_sc_hd__a21bo_1 c410 (.A1(clknet_1_0__leaf_net401),
    .A2(net291),
    .B1_N(net299),
    .X(net421));
 sky130_fd_sc_hd__xnor2_2 c411 (.A(net396),
    .B(net837),
    .Y(net422));
 sky130_fd_sc_hd__dfsbp_2 c412 (.CLK(clknet_leaf_2_clk),
    .D(clknet_1_1__leaf_net293),
    .SET_B(net414),
    .Q(net424),
    .Q_N(net423));
 sky130_fd_sc_hd__sdfxbp_1 c413 (.CLK(clknet_leaf_3_clk),
    .D(net415),
    .SCD(clknet_1_1__leaf_net421),
    .SCE(net423),
    .Q(net426),
    .Q_N(net425));
 sky130_fd_sc_hd__sdfxtp_1 c414 (.CLK(clknet_leaf_34_clk),
    .D(net418),
    .SCD(net414),
    .SCE(net909),
    .Q(net427));
 sky130_fd_sc_hd__sdfxtp_2 c415 (.CLK(clknet_leaf_3_clk),
    .D(net391),
    .SCD(net420),
    .SCE(net423),
    .Q(net428));
 sky130_fd_sc_hd__a21bo_1 c416 (.A1(net409),
    .A2(net420),
    .B1_N(net428),
    .X(net429));
 sky130_fd_sc_hd__mux4_1 c417 (.A0(clknet_1_0__leaf_net421),
    .A1(net273),
    .A2(net409),
    .A3(net411),
    .S0(net290),
    .S1(net414),
    .X(net430));
 sky130_fd_sc_hd__mux4_1 c418 (.A0(net425),
    .A1(net429),
    .A2(net297),
    .A3(net411),
    .S0(net414),
    .S1(net766),
    .X(net431));
 sky130_fd_sc_hd__sdfxtp_1 c419 (.CLK(clknet_leaf_2_clk),
    .D(net12),
    .SCD(net766),
    .SCE(net767),
    .Q(net432));
 sky130_fd_sc_hd__buf_1 c42 (.A(net41),
    .X(net18));
 sky130_fd_sc_hd__buf_1 c420 (.A(net753),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_1 c421 (.A(net753),
    .X(net434));
 sky130_fd_sc_hd__xnor2_1 c422 (.A(clknet_1_0__leaf_net303),
    .B(net411),
    .Y(net435));
 sky130_fd_sc_hd__xnor2_2 c423 (.A(net433),
    .B(net36),
    .Y(net436));
 sky130_fd_sc_hd__xnor2_2 c424 (.A(net416),
    .B(net423),
    .Y(net437));
 sky130_fd_sc_hd__dfbbn_1 c425 (.CLK_N(clknet_leaf_1_clk),
    .D(net166),
    .RESET_B(net436),
    .SET_B(net437),
    .Q(net438));
 sky130_fd_sc_hd__sdfrtp_1 c426 (.CLK(clknet_leaf_0_clk),
    .D(net856),
    .RESET_B(net12),
    .SCD(net411),
    .SCE(net393),
    .Q(net439));
 sky130_fd_sc_hd__dfstp_1 c427 (.CLK(clknet_leaf_1_clk),
    .D(net437),
    .SET_B(net805),
    .Q(net440));
 sky130_fd_sc_hd__xnor2_1 c428 (.A(net434),
    .B(net439),
    .Y(net441));
 sky130_fd_sc_hd__xnor2_1 c429 (.A(net439),
    .B(clknet_1_0__leaf_net435),
    .Y(net442));
 sky130_fd_sc_hd__xnor2_2 c43 (.A(net18),
    .B(net5),
    .Y(net19));
 sky130_fd_sc_hd__xnor2_1 c430 (.A(net441),
    .B(clknet_1_1__leaf_net303),
    .Y(net443));
 sky130_fd_sc_hd__dfstp_1 c431 (.CLK(clknet_leaf_1_clk),
    .D(net442),
    .SET_B(net899),
    .Q(net444));
 sky130_fd_sc_hd__a21bo_2 c432 (.A1(net412),
    .A2(net297),
    .B1_N(net393),
    .X(net445));
 sky130_fd_sc_hd__mux4_1 c433 (.A0(clknet_1_1__leaf_net435),
    .A1(net444),
    .A2(net445),
    .A3(net252),
    .S0(net312),
    .S1(net437),
    .X(net446));
 sky130_fd_sc_hd__mux4_1 c434 (.A0(net444),
    .A1(net437),
    .A2(net322),
    .A3(net252),
    .S0(net436),
    .S1(net768),
    .X(net447));
 sky130_fd_sc_hd__a21bo_1 c435 (.A1(clknet_1_1__leaf_net443),
    .A2(net444),
    .B1_N(net768),
    .X(net448));
 sky130_fd_sc_hd__xnor2_1 c436 (.A(net436),
    .B(net444),
    .Y(net449));
 sky130_fd_sc_hd__sdfrtp_1 c437 (.CLK(clknet_leaf_1_clk),
    .D(net449),
    .RESET_B(net859),
    .SCD(clknet_1_0__leaf_net448),
    .SCE(net968),
    .Q(net450));
 sky130_fd_sc_hd__xnor2_1 c438 (.A(net438),
    .B(clknet_1_0__leaf_net443),
    .Y(net451));
 sky130_fd_sc_hd__dfstp_4 c439 (.CLK(clknet_leaf_1_clk),
    .D(net449),
    .SET_B(net851),
    .Q(net816));
 sky130_fd_sc_hd__dfrbp_1 c44 (.CLK(clknet_leaf_31_clk),
    .D(net33),
    .RESET_B(net844),
    .Q(net21),
    .Q_N(net20));
 sky130_fd_sc_hd__mux4_1 c440 (.A0(net394),
    .A1(clknet_1_0__leaf_net451),
    .A2(net816),
    .A3(net414),
    .S0(net444),
    .S1(net769),
    .X(net452));
 sky130_fd_sc_hd__a21bo_1 c441 (.A1(net186),
    .A2(net424),
    .B1_N(net34),
    .X(net453));
 sky130_fd_sc_hd__dfbbn_1 c442 (.CLK_N(clknet_leaf_1_clk),
    .D(net318),
    .RESET_B(net407),
    .SET_B(net920),
    .Q(net455),
    .Q_N(net454));
 sky130_fd_sc_hd__buf_1 c443 (.A(net746),
    .X(net456));
 sky130_fd_sc_hd__dfbbp_1 c444 (.CLK(clknet_leaf_12_clk),
    .D(net327),
    .RESET_B(net456),
    .SET_B(clknet_1_1__leaf_net294),
    .Q(net458),
    .Q_N(net457));
 sky130_fd_sc_hd__a21bo_1 c445 (.A1(net408),
    .A2(net454),
    .B1_N(net339),
    .X(net459));
 sky130_fd_sc_hd__sdfxbp_1 c446 (.CLK(clknet_leaf_29_clk),
    .D(net877),
    .SCD(net459),
    .SCE(clknet_1_1__leaf_net187),
    .Q(net461),
    .Q_N(net460));
 sky130_fd_sc_hd__xnor2_1 c447 (.A(net461),
    .B(net769),
    .Y(net462));
 sky130_fd_sc_hd__buf_2 c448 (.A(net746),
    .X(net463));
 sky130_fd_sc_hd__sdfxbp_1 c449 (.CLK(clknet_leaf_1_clk),
    .D(clknet_1_1__leaf_net448),
    .SCD(net181),
    .SCE(net463),
    .Q(net465),
    .Q_N(net464));
 sky130_fd_sc_hd__clkbuf_4 c45 (.A(net39),
    .X(net22));
 sky130_fd_sc_hd__xnor2_1 c450 (.A(net312),
    .B(net463),
    .Y(net466));
 sky130_fd_sc_hd__a31o_1 c451 (.A1(net34),
    .A2(net436),
    .A3(net463),
    .B1(net462),
    .X(net467));
 sky130_fd_sc_hd__xnor2_1 c452 (.A(net36),
    .B(net464),
    .Y(net468));
 sky130_fd_sc_hd__a21bo_1 c453 (.A1(net465),
    .A2(net408),
    .B1_N(net463),
    .X(net469));
 sky130_fd_sc_hd__a31o_1 c454 (.A1(net27),
    .A2(net469),
    .A3(net466),
    .B1(net428),
    .X(net470));
 sky130_fd_sc_hd__a31o_1 c455 (.A1(net466),
    .A2(net345),
    .A3(net460),
    .B1(net463),
    .X(net471));
 sky130_fd_sc_hd__sdfxtp_1 c456 (.CLK(clknet_leaf_18_clk),
    .D(net470),
    .SCD(net471),
    .SCE(net468),
    .Q(net472));
 sky130_fd_sc_hd__sdfsbp_1 c457 (.CLK(clknet_leaf_18_clk),
    .D(net471),
    .SCD(net467),
    .SCE(net411),
    .SET_B(net414),
    .Q(net473));
 sky130_fd_sc_hd__sdfsbp_1 c458 (.CLK(clknet_leaf_18_clk),
    .D(net462),
    .SCD(net150),
    .SCE(net470),
    .SET_B(net905),
    .Q(net475),
    .Q_N(net474));
 sky130_fd_sc_hd__a21bo_1 c459 (.A1(net473),
    .A2(net463),
    .B1_N(net472),
    .X(net476));
 sky130_fd_sc_hd__dfbbn_2 c46 (.CLK_N(clknet_leaf_31_clk),
    .D(net18),
    .RESET_B(net38),
    .SET_B(net19),
    .Q(net24),
    .Q_N(net23));
 sky130_fd_sc_hd__sdfbbn_1 c460 (.CLK_N(clknet_leaf_12_clk),
    .D(net459),
    .RESET_B(net471),
    .SCD(net469),
    .SCE(net453),
    .SET_B(net191),
    .Q(net477));
 sky130_fd_sc_hd__a41o_1 c461 (.A1(net472),
    .A2(net337),
    .A3(net468),
    .A4(net463),
    .B1(net47),
    .X(net478));
 sky130_fd_sc_hd__a21bo_1 c462 (.A1(net298),
    .A2(net13),
    .B1_N(net476),
    .X(net479));
 sky130_fd_sc_hd__buf_1 c463 (.A(net740),
    .X(net817));
 sky130_fd_sc_hd__xnor2_2 c464 (.A(net339),
    .B(net860),
    .Y(net480));
 sky130_fd_sc_hd__xnor2_1 c465 (.A(net229),
    .B(net764),
    .Y(net481));
 sky130_fd_sc_hd__clkbuf_1 c466 (.A(net740),
    .X(net482));
 sky130_fd_sc_hd__dlrbn_1 c467 (.D(net455),
    .GATE_N(clknet_leaf_18_clk),
    .RESET_B(net480),
    .Q(net483));
 sky130_fd_sc_hd__xnor2_1 c468 (.A(net479),
    .B(net816),
    .Y(net484));
 sky130_fd_sc_hd__dlrbn_1 c469 (.D(net468),
    .GATE_N(clknet_leaf_18_clk),
    .RESET_B(net356),
    .Q(net485));
 sky130_fd_sc_hd__xnor2_4 c47 (.A(net24),
    .B(net928),
    .Y(net25));
 sky130_fd_sc_hd__dlrbp_1 c470 (.D(net476),
    .GATE(clknet_leaf_20_clk),
    .RESET_B(net484),
    .Q(net486));
 sky130_fd_sc_hd__xnor2_2 c471 (.A(net344),
    .B(net835),
    .Y(net487));
 sky130_fd_sc_hd__xnor2_2 c472 (.A(net485),
    .B(net298),
    .Y(net488));
 sky130_fd_sc_hd__dlrbp_1 c473 (.D(net487),
    .GATE(clknet_leaf_18_clk),
    .RESET_B(net362),
    .Q(net489));
 sky130_fd_sc_hd__xnor2_1 c474 (.A(net863),
    .B(net455),
    .Y(net490));
 sky130_fd_sc_hd__sdfxtp_2 c475 (.CLK(clknet_leaf_17_clk),
    .D(net207),
    .SCD(net251),
    .SCE(net467),
    .Q(net491));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(net388),
    .A1(net207),
    .A2(net414),
    .A3(net488),
    .S0(net362),
    .S1(net480),
    .X(net492));
 sky130_fd_sc_hd__sdfxtp_1 c477 (.CLK(clknet_leaf_19_clk),
    .D(net140),
    .SCD(net360),
    .SCE(net896),
    .Q(net493));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(net480),
    .A1(net251),
    .A2(net490),
    .A3(net360),
    .S0(net952),
    .S1(net967),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(net478),
    .A1(net487),
    .A2(net491),
    .A3(net835),
    .S0(net388),
    .S1(net54),
    .X(net495));
 sky130_fd_sc_hd__dfrbp_2 c48 (.CLK(clknet_leaf_26_clk),
    .D(net19),
    .RESET_B(net850),
    .Q(net832),
    .Q_N(net26));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net943),
    .A1(net480),
    .A2(net207),
    .A3(net487),
    .S0(net360),
    .S1(net966),
    .X(net496));
 sky130_fd_sc_hd__a21bo_1 c481 (.A1(net483),
    .A2(net481),
    .B1_N(net47),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(net150),
    .A1(net497),
    .A2(net487),
    .A3(net484),
    .S0(net773),
    .S1(net775),
    .X(net498));
 sky130_fd_sc_hd__a21bo_1 c487 (.A1(net406),
    .A2(net385),
    .B1_N(net491),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_1 c488 (.A(net784),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_1 c489 (.A(net784),
    .X(net818));
 sky130_fd_sc_hd__xnor2_4 c49 (.A(net30),
    .B(net25),
    .Y(net27));
 sky130_fd_sc_hd__a21bo_1 c490 (.A1(net499),
    .A2(net500),
    .B1_N(net840),
    .X(net501));
 sky130_fd_sc_hd__dfbbn_1 c491 (.CLK_N(clknet_leaf_21_clk),
    .D(clknet_1_1__leaf_net233),
    .RESET_B(net493),
    .SET_B(clknet_1_0__leaf_net827),
    .Q(net810));
 sky130_fd_sc_hd__dfbbn_1 c492 (.CLK_N(clknet_leaf_16_clk),
    .D(net501),
    .RESET_B(net816),
    .SET_B(clknet_1_1__leaf_net372),
    .Q(net822));
 sky130_fd_sc_hd__dfbbp_1 c493 (.CLK(clknet_leaf_20_clk),
    .D(net92),
    .RESET_B(net841),
    .SET_B(clknet_1_0__leaf_net372),
    .Q(net502));
 sky130_fd_sc_hd__sdfxbp_1 c494 (.CLK(clknet_leaf_20_clk),
    .D(net378),
    .SCD(net834),
    .SCE(net841),
    .Q(net504),
    .Q_N(net503));
 sky130_fd_sc_hd__a41o_1 c495 (.A1(net373),
    .A2(net491),
    .A3(net432),
    .A4(net503),
    .B1(net217),
    .X(net505));
 sky130_fd_sc_hd__sdfxbp_1 c496 (.CLK(clknet_leaf_16_clk),
    .D(net841),
    .SCD(net432),
    .SCE(clknet_1_1__leaf_net372),
    .Q(net826));
 sky130_fd_sc_hd__a21bo_1 c497 (.A1(net486),
    .A2(net236),
    .B1_N(net504),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(net502),
    .A1(net151),
    .A2(net406),
    .A3(net823),
    .S0(net503),
    .S1(net384),
    .X(net507));
 sky130_fd_sc_hd__sdfxtp_1 c499 (.CLK(clknet_leaf_19_clk),
    .D(net414),
    .SCD(net813),
    .SCE(net829),
    .Q(net508));
 sky130_fd_sc_hd__xnor2_4 c50 (.A(net25),
    .B(net22),
    .Y(net28));
 sky130_fd_sc_hd__a21bo_1 c500 (.A1(net505),
    .A2(net367),
    .B1_N(net504),
    .X(net509));
 sky130_fd_sc_hd__sdfxtp_1 c501 (.CLK(clknet_leaf_19_clk),
    .D(net356),
    .SCD(net892),
    .SCE(net834),
    .Q(net824));
 sky130_fd_sc_hd__a21bo_1 c502 (.A1(net506),
    .A2(net504),
    .B1_N(net491),
    .X(net825));
 sky130_fd_sc_hd__sdfbbp_1 c503 (.CLK(clknet_leaf_16_clk),
    .D(net432),
    .RESET_B(net509),
    .SCD(net257),
    .SCE(net503),
    .SET_B(net816));
 sky130_fd_sc_hd__clkbuf_2 c504 (.A(net737),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_4 c505 (.A(net737),
    .X(net511));
 sky130_fd_sc_hd__xnor2_1 c506 (.A(net793),
    .B(net511),
    .Y(net512));
 sky130_fd_sc_hd__buf_1 c507 (.A(net124),
    .X(net513));
 sky130_fd_sc_hd__clkbuf_1 c508 (.A(net836),
    .X(net514));
 sky130_fd_sc_hd__buf_2 c509 (.A(net802),
    .X(net515));
 sky130_fd_sc_hd__xnor2_2 c51 (.A(net22),
    .B(net27),
    .Y(net29));
 sky130_fd_sc_hd__xnor2_4 c510 (.A(net121),
    .B(net402),
    .Y(net516));
 sky130_fd_sc_hd__xnor2_1 c511 (.A(net402),
    .B(net793),
    .Y(net517));
 sky130_fd_sc_hd__xnor2_1 c512 (.A(clknet_1_1__leaf_net267),
    .B(net515),
    .Y(net518));
 sky130_fd_sc_hd__clkbuf_1 c513 (.A(net386),
    .X(net519));
 sky130_fd_sc_hd__clkbuf_2 c514 (.A(net785),
    .X(net520));
 sky130_fd_sc_hd__xnor2_1 c515 (.A(net518),
    .B(net520),
    .Y(net521));
 sky130_fd_sc_hd__dlrtn_1 c516 (.D(net519),
    .GATE_N(clknet_leaf_4_clk),
    .RESET_B(net520),
    .Q(net522));
 sky130_fd_sc_hd__xnor2_1 c517 (.A(net520),
    .B(net387),
    .Y(net523));
 sky130_fd_sc_hd__dlrtn_2 c518 (.D(net523),
    .GATE_N(clknet_leaf_4_clk),
    .RESET_B(net512),
    .Q(net524));
 sky130_fd_sc_hd__dlrtn_4 c519 (.D(net522),
    .GATE_N(clknet_leaf_5_clk),
    .RESET_B(net513),
    .Q(net525));
 sky130_fd_sc_hd__buf_2 c52 (.A(net794),
    .X(net30));
 sky130_fd_sc_hd__xnor2_1 c520 (.A(net517),
    .B(net525),
    .Y(net526));
 sky130_fd_sc_hd__xnor2_1 c521 (.A(net525),
    .B(net911),
    .Y(net527));
 sky130_fd_sc_hd__xnor2_1 c522 (.A(net512),
    .B(net520),
    .Y(net528));
 sky130_fd_sc_hd__dlrtp_1 c523 (.D(net514),
    .GATE(clknet_leaf_5_clk),
    .RESET_B(net527),
    .Q(net529));
 sky130_fd_sc_hd__xnor2_1 c524 (.A(net528),
    .B(net387),
    .Y(net530));
 sky130_fd_sc_hd__buf_1 c525 (.A(clknet_1_1__leaf_net139),
    .X(net531));
 sky130_fd_sc_hd__clkbuf_2 c526 (.A(net745),
    .X(net532));
 sky130_fd_sc_hd__sdfxtp_1 c527 (.CLK(clknet_leaf_2_clk),
    .D(net531),
    .SCD(net395),
    .SCE(clknet_1_0__leaf_net279),
    .Q(net533));
 sky130_fd_sc_hd__xnor2_1 c528 (.A(net964),
    .B(net428),
    .Y(net534));
 sky130_fd_sc_hd__xnor2_1 c529 (.A(clknet_1_1__leaf_net142),
    .B(net524),
    .Y(net535));
 sky130_fd_sc_hd__buf_2 c53 (.A(net789),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 c530 (.A(net744),
    .X(net536));
 sky130_fd_sc_hd__xnor2_1 c531 (.A(net536),
    .B(net427),
    .Y(net537));
 sky130_fd_sc_hd__xnor2_2 c532 (.A(net276),
    .B(net536),
    .Y(net538));
 sky130_fd_sc_hd__a21bo_1 c533 (.A1(net536),
    .A2(net532),
    .B1_N(net422),
    .X(net539));
 sky130_fd_sc_hd__dlrtp_2 c534 (.D(net514),
    .GATE(clknet_leaf_5_clk),
    .RESET_B(net395),
    .Q(net540));
 sky130_fd_sc_hd__dlrtp_1 c535 (.D(clknet_1_1__leaf_net279),
    .GATE(clknet_leaf_2_clk),
    .RESET_B(clknet_1_0__leaf_net535),
    .Q(net541));
 sky130_fd_sc_hd__edfxbp_1 c536 (.CLK(clknet_leaf_5_clk),
    .D(net513),
    .DE(net539),
    .Q(net543),
    .Q_N(net542));
 sky130_fd_sc_hd__xnor2_1 c537 (.A(net526),
    .B(net135),
    .Y(net544));
 sky130_fd_sc_hd__a21bo_1 c538 (.A1(net300),
    .A2(net536),
    .B1_N(net273),
    .X(net545));
 sky130_fd_sc_hd__a21bo_1 c539 (.A1(net538),
    .A2(net422),
    .B1_N(net543),
    .X(net546));
 sky130_fd_sc_hd__a21bo_1 c54 (.A1(net11),
    .A2(net798),
    .B1_N(net15),
    .X(net32));
 sky130_fd_sc_hd__dfbbn_2 c540 (.CLK_N(clknet_leaf_2_clk),
    .D(net539),
    .RESET_B(net395),
    .SET_B(net513),
    .Q(net548),
    .Q_N(net547));
 sky130_fd_sc_hd__edfxtp_1 c541 (.CLK(clknet_leaf_5_clk),
    .D(net544),
    .DE(net542),
    .Q(net549));
 sky130_fd_sc_hd__xnor2_1 c542 (.A(net422),
    .B(net397),
    .Y(net828));
 sky130_fd_sc_hd__mux4_1 c543 (.A0(net803),
    .A1(net539),
    .A2(net828),
    .A3(net545),
    .S0(net544),
    .S1(net540),
    .X(net550));
 sky130_fd_sc_hd__dfbbn_1 c544 (.CLK_N(clknet_leaf_5_clk),
    .D(net427),
    .RESET_B(net549),
    .SET_B(net544),
    .Q(net552),
    .Q_N(net551));
 sky130_fd_sc_hd__dfbbp_1 c545 (.CLK(clknet_leaf_2_clk),
    .D(net395),
    .RESET_B(net552),
    .SET_B(net539),
    .Q(net554),
    .Q_N(net553));
 sky130_fd_sc_hd__xnor2_4 c546 (.A(net445),
    .B(net424),
    .Y(net555));
 sky130_fd_sc_hd__sdlclkp_1 c547 (.CLK(clknet_leaf_12_clk),
    .GATE(net266),
    .SCE(net29),
    .GCLK(net556));
 sky130_fd_sc_hd__sdfstp_1 c548 (.CLK(clknet_leaf_2_clk),
    .D(net787),
    .SCD(net915),
    .SCE(clknet_1_0__leaf_net287),
    .SET_B(net252),
    .Q(net557));
 sky130_fd_sc_hd__xnor2_4 c549 (.A(net861),
    .B(net547),
    .Y(net558));
 sky130_fd_sc_hd__clkbuf_1 c55 (.A(net32),
    .X(net33));
 sky130_fd_sc_hd__sdlclkp_2 c550 (.CLK(clknet_leaf_11_clk),
    .GATE(clknet_1_0__leaf_net521),
    .SCE(net914),
    .GCLK(net559));
 sky130_fd_sc_hd__xnor2_1 c551 (.A(net816),
    .B(net777),
    .Y(net560));
 sky130_fd_sc_hd__sdlclkp_4 c552 (.CLK(clknet_leaf_11_clk),
    .GATE(net151),
    .SCE(net555),
    .GCLK(net561));
 sky130_fd_sc_hd__xnor2_1 c553 (.A(net555),
    .B(net524),
    .Y(net562));
 sky130_fd_sc_hd__xnor2_2 c554 (.A(net554),
    .B(net540),
    .Y(net563));
 sky130_fd_sc_hd__dfrbp_1 c555 (.CLK(clknet_leaf_12_clk),
    .D(net29),
    .RESET_B(net307),
    .Q(net564));
 sky130_fd_sc_hd__dfrbp_1 c556 (.CLK(clknet_leaf_9_clk),
    .D(net563),
    .RESET_B(net813),
    .Q(net821),
    .Q_N(net565));
 sky130_fd_sc_hd__dfrtn_1 c557 (.CLK_N(clknet_leaf_2_clk),
    .D(clknet_1_1__leaf_net451),
    .RESET_B(net428),
    .Q(net566));
 sky130_fd_sc_hd__sdfbbn_1 c558 (.CLK_N(clknet_leaf_2_clk),
    .D(net560),
    .RESET_B(clknet_1_0__leaf_net294),
    .SCD(net563),
    .SCE(net524),
    .SET_B(net510),
    .Q(net568),
    .Q_N(net567));
 sky130_fd_sc_hd__dfrtp_1 c559 (.CLK(clknet_leaf_11_clk),
    .D(net252),
    .RESET_B(net307),
    .Q(net569));
 sky130_fd_sc_hd__dfrtn_1 c56 (.CLK_N(clknet_leaf_31_clk),
    .D(net30),
    .RESET_B(net0),
    .Q(net34));
 sky130_fd_sc_hd__a41o_1 c560 (.A1(net273),
    .A2(net923),
    .A3(net555),
    .A4(net565),
    .B1(net558),
    .X(net570));
 sky130_fd_sc_hd__mux4_1 c561 (.A0(net853),
    .A1(net568),
    .A2(net563),
    .A3(net532),
    .S0(net555),
    .S1(net157),
    .X(net571));
 sky130_fd_sc_hd__xnor2_1 c562 (.A(net564),
    .B(net313),
    .Y(net572));
 sky130_fd_sc_hd__a21bo_1 c563 (.A1(net306),
    .A2(net816),
    .B1_N(net771),
    .X(net573));
 sky130_fd_sc_hd__sdfbbn_1 c564 (.CLK_N(clknet_leaf_11_clk),
    .D(net450),
    .RESET_B(net570),
    .SCD(net563),
    .SCE(net566),
    .SET_B(net555),
    .Q(net575),
    .Q_N(net574));
 sky130_fd_sc_hd__dfrtp_1 c565 (.CLK(clknet_leaf_11_clk),
    .D(net163),
    .RESET_B(net854),
    .Q(net576));
 sky130_fd_sc_hd__sdfbbp_1 c566 (.CLK(clknet_leaf_11_clk),
    .D(net890),
    .RESET_B(net555),
    .SCD(net567),
    .SCE(net524),
    .SET_B(clknet_1_1__leaf_net521),
    .Q(net578),
    .Q_N(net577));
 sky130_fd_sc_hd__xnor2_1 c567 (.A(net203),
    .B(net541),
    .Y(net579));
 sky130_fd_sc_hd__clkbuf_1 c568 (.A(net743),
    .X(net580));
 sky130_fd_sc_hd__a21bo_1 c569 (.A1(net580),
    .A2(net857),
    .B1_N(net572),
    .X(net581));
 sky130_fd_sc_hd__buf_1 c57 (.A(net32),
    .X(net35));
 sky130_fd_sc_hd__a21bo_1 c570 (.A1(net869),
    .A2(net397),
    .B1_N(net834),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_1 c571 (.A(net954),
    .X(net583));
 sky130_fd_sc_hd__a21bo_1 c572 (.A1(net556),
    .A2(clknet_1_1__leaf_net287),
    .B1_N(net816),
    .X(net584));
 sky130_fd_sc_hd__sdfxbp_1 c573 (.CLK(clknet_leaf_12_clk),
    .D(net314),
    .SCD(net135),
    .SCE(clknet_1_1__leaf_net202),
    .Q(net585));
 sky130_fd_sc_hd__a21bo_1 c574 (.A1(net461),
    .A2(net835),
    .B1_N(net816),
    .X(net586));
 sky130_fd_sc_hd__xnor2_1 c575 (.A(clknet_1_1__leaf_net287),
    .B(net203),
    .Y(net587));
 sky130_fd_sc_hd__xnor2_1 c576 (.A(net458),
    .B(net511),
    .Y(net588));
 sky130_fd_sc_hd__sdfxbp_1 c577 (.CLK(clknet_leaf_18_clk),
    .D(net47),
    .SCD(net587),
    .SCE(net586),
    .Q(net589));
 sky130_fd_sc_hd__sdfxtp_1 c578 (.CLK(clknet_leaf_13_clk),
    .D(net583),
    .SCD(net582),
    .SCE(net586),
    .Q(net590));
 sky130_fd_sc_hd__dfrtp_1 c579 (.CLK(clknet_leaf_12_clk),
    .D(net874),
    .RESET_B(net870),
    .Q(net591));
 sky130_fd_sc_hd__xnor2_4 c58 (.A(net804),
    .B(net801),
    .Y(net36));
 sky130_fd_sc_hd__xnor2_1 c580 (.A(net579),
    .B(net307),
    .Y(net592));
 sky130_fd_sc_hd__xnor2_2 c581 (.A(net589),
    .B(net762),
    .Y(net593));
 sky130_fd_sc_hd__sdfxtp_1 c582 (.CLK(clknet_leaf_12_clk),
    .D(net884),
    .SCD(net938),
    .SCE(net545),
    .Q(net594));
 sky130_fd_sc_hd__a41o_1 c583 (.A1(net586),
    .A2(net946),
    .A3(net816),
    .A4(net591),
    .B1(net510),
    .X(net595));
 sky130_fd_sc_hd__sdfxtp_1 c584 (.CLK(clknet_leaf_12_clk),
    .D(net595),
    .SCD(net588),
    .SCE(net925),
    .Q(net596));
 sky130_fd_sc_hd__dfbbn_1 c585 (.CLK_N(clknet_leaf_11_clk),
    .D(net533),
    .RESET_B(net572),
    .SET_B(clknet_1_1__leaf_net294),
    .Q(net598),
    .Q_N(net597));
 sky130_fd_sc_hd__a41o_1 c586 (.A1(net598),
    .A2(net596),
    .A3(net457),
    .A4(net594),
    .B1(clknet_1_1__leaf_net287),
    .X(net599));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(net545),
    .A1(net599),
    .A2(net597),
    .A3(net586),
    .S0(net591),
    .S1(net593),
    .X(net600));
 sky130_fd_sc_hd__dfbbn_1 c588 (.CLK_N(clknet_leaf_17_clk),
    .D(net482),
    .RESET_B(net69),
    .SET_B(net775),
    .Q(net601));
 sky130_fd_sc_hd__xnor2_1 c589 (.A(net559),
    .B(net601),
    .Y(net602));
 sky130_fd_sc_hd__xnor2_1 c59 (.A(net31),
    .B(net15),
    .Y(net37));
 sky130_fd_sc_hd__sdfbbn_1 c590 (.CLK_N(clknet_leaf_17_clk),
    .D(net365),
    .RESET_B(net602),
    .SCD(net217),
    .SCE(net69),
    .SET_B(net832),
    .Q(net603));
 sky130_fd_sc_hd__a21bo_1 c591 (.A1(net510),
    .A2(net477),
    .B1_N(net775),
    .X(net604));
 sky130_fd_sc_hd__xnor2_1 c592 (.A(net428),
    .B(net578),
    .Y(net605));
 sky130_fd_sc_hd__buf_1 c593 (.A(net965),
    .X(net606));
 sky130_fd_sc_hd__clkbuf_1 c594 (.A(net924),
    .X(net607));
 sky130_fd_sc_hd__dfbbp_1 c595 (.CLK(clknet_leaf_17_clk),
    .D(net582),
    .RESET_B(clknet_1_1__leaf_net187),
    .SET_B(net775),
    .Q(net608));
 sky130_fd_sc_hd__xnor2_1 c596 (.A(net524),
    .B(net605),
    .Y(net609));
 sky130_fd_sc_hd__sdfxbp_1 c597 (.CLK(clknet_leaf_12_clk),
    .D(net912),
    .SCD(net117),
    .SCE(net360),
    .Q(net610));
 sky130_fd_sc_hd__a21bo_1 c598 (.A1(net789),
    .A2(net603),
    .B1_N(net834),
    .X(net611));
 sky130_fd_sc_hd__a21bo_1 c599 (.A1(net540),
    .A2(net609),
    .B1_N(net397),
    .X(net831));
 sky130_fd_sc_hd__dfxbp_1 c60 (.CLK(clknet_leaf_25_clk),
    .D(net35),
    .Q(net39),
    .Q_N(net38));
 sky130_fd_sc_hd__sdfxbp_1 c600 (.CLK(clknet_leaf_17_clk),
    .D(net611),
    .SCD(net607),
    .SCE(net251),
    .Q(net612));
 sky130_fd_sc_hd__a21bo_1 c601 (.A1(net610),
    .A2(net612),
    .B1_N(net540),
    .X(net613));
 sky130_fd_sc_hd__sdfbbn_1 c602 (.CLK_N(clknet_leaf_17_clk),
    .D(net219),
    .RESET_B(net608),
    .SCD(net488),
    .SCE(net606),
    .SET_B(net69),
    .Q(net614));
 sky130_fd_sc_hd__a21bo_1 c603 (.A1(net930),
    .A2(net613),
    .B1_N(net787),
    .X(net615));
 sky130_fd_sc_hd__sdfxtp_1 c604 (.CLK(clknet_leaf_13_clk),
    .D(net592),
    .SCD(net615),
    .SCE(net497),
    .Q(net616));
 sky130_fd_sc_hd__sdfxtp_1 c605 (.CLK(clknet_leaf_17_clk),
    .D(clknet_1_1__leaf_net187),
    .SCD(net497),
    .SCE(net362),
    .Q(net617));
 sky130_fd_sc_hd__sdfxtp_1 c606 (.CLK(clknet_leaf_17_clk),
    .D(clknet_1_1__leaf_net202),
    .SCD(net958),
    .SCE(net614),
    .Q(net618));
 sky130_fd_sc_hd__xnor2_1 c607 (.A(net618),
    .B(net617),
    .Y(net619));
 sky130_fd_sc_hd__a21bo_1 c608 (.A1(net619),
    .A2(net548),
    .B1_N(net616),
    .X(net620));
 sky130_fd_sc_hd__clkbuf_1 c61 (.A(net34),
    .X(net40));
 sky130_fd_sc_hd__dfrtp_4 c62 (.CLK(clknet_leaf_31_clk),
    .D(net33),
    .RESET_B(net30),
    .Q(net41));
 sky130_fd_sc_hd__buf_1 c63 (.A(net21),
    .X(net42));
 sky130_fd_sc_hd__xnor2_4 c630 (.A(net266),
    .B(net525),
    .Y(net621));
 sky130_fd_sc_hd__clkbuf_1 c631 (.A(net517),
    .X(net622));
 sky130_fd_sc_hd__clkbuf_1 c632 (.A(net621),
    .X(net623));
 sky130_fd_sc_hd__xnor2_1 c633 (.A(net387),
    .B(net621),
    .Y(net624));
 sky130_fd_sc_hd__xnor2_2 c634 (.A(net621),
    .B(net118),
    .Y(net625));
 sky130_fd_sc_hd__xnor2_4 c635 (.A(net525),
    .B(net397),
    .Y(net626));
 sky130_fd_sc_hd__xnor2_1 c636 (.A(net263),
    .B(net626),
    .Y(net627));
 sky130_fd_sc_hd__dfsbp_1 c637 (.CLK(clknet_leaf_5_clk),
    .D(net530),
    .SET_B(net253),
    .Q(net628));
 sky130_fd_sc_hd__dfbbn_1 c638 (.CLK_N(clknet_leaf_5_clk),
    .D(net623),
    .RESET_B(net118),
    .SET_B(net263),
    .Q(net629));
 sky130_fd_sc_hd__clkbuf_1 c639 (.A(net527),
    .X(net630));
 sky130_fd_sc_hd__clkbuf_4 c64 (.A(net25),
    .X(net43));
 sky130_fd_sc_hd__xnor2_4 c640 (.A(net796),
    .B(net621),
    .Y(net631));
 sky130_fd_sc_hd__dfsbp_2 c641 (.CLK(clknet_leaf_6_clk),
    .D(net627),
    .SET_B(net631),
    .Q(net633),
    .Q_N(net632));
 sky130_fd_sc_hd__xnor2_1 c642 (.A(net630),
    .B(net118),
    .Y(net634));
 sky130_fd_sc_hd__dfstp_1 c643 (.CLK(clknet_leaf_6_clk),
    .D(net253),
    .SET_B(net626),
    .Q(net635));
 sky130_fd_sc_hd__dfstp_1 c644 (.CLK(clknet_leaf_7_clk),
    .D(net631),
    .SET_B(net855),
    .Q(net636));
 sky130_fd_sc_hd__xnor2_1 c645 (.A(net951),
    .B(net837),
    .Y(net637));
 sky130_fd_sc_hd__a21bo_1 c646 (.A1(net622),
    .A2(net266),
    .B1_N(net632),
    .X(net638));
 sky130_fd_sc_hd__a21bo_1 c647 (.A1(net947),
    .A2(net525),
    .B1_N(net621),
    .X(net639));
 sky130_fd_sc_hd__dfstp_1 c648 (.CLK(clknet_leaf_6_clk),
    .D(net639),
    .SET_B(net638),
    .Q(net640));
 sky130_fd_sc_hd__sdfstp_1 c649 (.CLK(clknet_leaf_5_clk),
    .D(net404),
    .SCD(net633),
    .SCE(net638),
    .SET_B(net387),
    .Q(net641));
 sky130_fd_sc_hd__mux4_1 c65 (.A0(net65),
    .A1(net58),
    .A2(net64),
    .A3(net43),
    .S0(net31),
    .S1(clknet_1_0__leaf_net757),
    .X(net44));
 sky130_fd_sc_hd__dfbbn_2 c650 (.CLK_N(clknet_leaf_5_clk),
    .D(net637),
    .RESET_B(net641),
    .SET_B(net253),
    .Q(net643),
    .Q_N(net642));
 sky130_fd_sc_hd__dlrbn_1 c651 (.D(net546),
    .GATE_N(clknet_leaf_7_clk),
    .RESET_B(net515),
    .Q(net644));
 sky130_fd_sc_hd__xnor2_4 c652 (.A(net626),
    .B(net543),
    .Y(net645));
 sky130_fd_sc_hd__dlrbn_1 c653 (.D(net624),
    .GATE_N(clknet_leaf_6_clk),
    .RESET_B(net645),
    .Q(net646));
 sky130_fd_sc_hd__mux4_1 c654 (.A0(net640),
    .A1(net646),
    .A2(net551),
    .A3(net135),
    .S0(net546),
    .S1(net516),
    .X(net647));
 sky130_fd_sc_hd__dlrbp_1 c655 (.D(net543),
    .GATE(clknet_leaf_5_clk),
    .RESET_B(net546),
    .Q(net649),
    .Q_N(net648));
 sky130_fd_sc_hd__dfbbp_1 c656 (.CLK(clknet_leaf_7_clk),
    .D(net644),
    .RESET_B(net511),
    .SET_B(net645),
    .Q(net650));
 sky130_fd_sc_hd__sdfxbp_1 c657 (.CLK(clknet_leaf_7_clk),
    .D(net537),
    .SCD(net638),
    .SCE(net511),
    .Q(net652),
    .Q_N(net651));
 sky130_fd_sc_hd__xnor2_2 c658 (.A(net796),
    .B(net779),
    .Y(net653));
 sky130_fd_sc_hd__xnor2_1 c659 (.A(net552),
    .B(net626),
    .Y(net654));
 sky130_fd_sc_hd__dfbbp_1 c66 (.CLK(clknet_leaf_25_clk),
    .D(net44),
    .RESET_B(net42),
    .SET_B(net58),
    .Q(net46),
    .Q_N(net45));
 sky130_fd_sc_hd__a31o_1 c660 (.A1(net636),
    .A2(net652),
    .A3(net648),
    .B1(net113),
    .X(net655));
 sky130_fd_sc_hd__a21bo_1 c661 (.A1(net796),
    .A2(net649),
    .B1_N(net542),
    .X(net656));
 sky130_fd_sc_hd__xnor2_1 c662 (.A(net538),
    .B(net529),
    .Y(net657));
 sky130_fd_sc_hd__xnor2_1 c663 (.A(net529),
    .B(net651),
    .Y(net658));
 sky130_fd_sc_hd__sdfxbp_1 c664 (.CLK(clknet_leaf_7_clk),
    .D(net137),
    .SCD(net654),
    .SCE(net642),
    .Q(net659));
 sky130_fd_sc_hd__dlrbp_1 c665 (.D(net429),
    .GATE(clknet_leaf_7_clk),
    .RESET_B(net516),
    .Q(net661),
    .Q_N(net660));
 sky130_fd_sc_hd__xnor2_4 c666 (.A(net653),
    .B(net642),
    .Y(net662));
 sky130_fd_sc_hd__xnor2_1 c667 (.A(net957),
    .B(net662),
    .Y(net663));
 sky130_fd_sc_hd__xnor2_4 c668 (.A(net662),
    .B(net660),
    .Y(net664));
 sky130_fd_sc_hd__xnor2_1 c669 (.A(net652),
    .B(net756),
    .Y(net665));
 sky130_fd_sc_hd__xnor2_4 c67 (.A(net4),
    .B(net786),
    .Y(net47));
 sky130_fd_sc_hd__sdfxtp_1 c670 (.CLK(clknet_leaf_7_clk),
    .D(net956),
    .SCD(net944),
    .SCE(net664),
    .Q(net666));
 sky130_fd_sc_hd__dlrtn_1 c671 (.D(net665),
    .GATE_N(clknet_leaf_8_clk),
    .RESET_B(net645),
    .Q(net667));
 sky130_fd_sc_hd__buf_1 c672 (.A(net783),
    .X(net668));
 sky130_fd_sc_hd__sdfstp_1 c673 (.CLK(clknet_leaf_8_clk),
    .D(net634),
    .SCD(net668),
    .SCE(net651),
    .SET_B(net852),
    .Q(net669));
 sky130_fd_sc_hd__a21bo_1 c674 (.A1(net669),
    .A2(net668),
    .B1_N(net633),
    .X(net670));
 sky130_fd_sc_hd__clkbuf_1 c675 (.A(net783),
    .X(net671));
 sky130_fd_sc_hd__a21bo_1 c676 (.A1(net661),
    .A2(net670),
    .B1_N(net789),
    .X(net672));
 sky130_fd_sc_hd__sdfxtp_1 c677 (.CLK(clknet_leaf_8_clk),
    .D(net625),
    .SCD(net657),
    .SCE(net852),
    .Q(net673));
 sky130_fd_sc_hd__sdfxtp_1 c678 (.CLK(clknet_leaf_9_clk),
    .D(net658),
    .SCD(net135),
    .SCE(clknet_1_1__leaf_net535),
    .Q(net674));
 sky130_fd_sc_hd__sdfbbp_1 c679 (.CLK(clknet_leaf_9_clk),
    .D(net515),
    .RESET_B(net663),
    .SCD(net668),
    .SCE(net671),
    .SET_B(net864),
    .Q(net676),
    .Q_N(net675));
 sky130_fd_sc_hd__buf_1 c68 (.A(net42),
    .X(net48));
 sky130_fd_sc_hd__a21bo_1 c680 (.A1(net652),
    .A2(net657),
    .B1_N(net257),
    .X(net677));
 sky130_fd_sc_hd__a41o_1 c681 (.A1(net118),
    .A2(net643),
    .A3(net532),
    .A4(net515),
    .B1(net135),
    .X(net678));
 sky130_fd_sc_hd__dfbbn_1 c682 (.CLK_N(clknet_leaf_9_clk),
    .D(net638),
    .RESET_B(net645),
    .SET_B(net672),
    .Q(net679));
 sky130_fd_sc_hd__dfbbn_1 c683 (.CLK_N(clknet_leaf_7_clk),
    .D(net645),
    .RESET_B(net937),
    .SET_B(net677),
    .Q(net680));
 sky130_fd_sc_hd__dfbbp_1 c684 (.CLK(clknet_leaf_10_clk),
    .D(net655),
    .RESET_B(net664),
    .SET_B(net864),
    .Q(net682),
    .Q_N(net681));
 sky130_fd_sc_hd__sdfxbp_1 c685 (.CLK(clknet_leaf_10_clk),
    .D(net643),
    .SCD(net663),
    .SCE(net180),
    .Q(net683));
 sky130_fd_sc_hd__sdfxbp_1 c686 (.CLK(clknet_leaf_9_clk),
    .D(net410),
    .SCD(net664),
    .SCE(net682),
    .Q(net684));
 sky130_fd_sc_hd__a21bo_1 c687 (.A1(net678),
    .A2(net913),
    .B1_N(net515),
    .X(net685));
 sky130_fd_sc_hd__sdfbbn_1 c688 (.CLK_N(clknet_leaf_9_clk),
    .D(net936),
    .RESET_B(net799),
    .SCD(net516),
    .SCE(net674),
    .SET_B(net625),
    .Q(net687),
    .Q_N(net686));
 sky130_fd_sc_hd__sedfxbp_1 c689 (.CLK(clknet_leaf_9_clk),
    .D(net941),
    .DE(net684),
    .SCD(net927),
    .SCE(net677),
    .Q(net689),
    .Q_N(net688));
 sky130_fd_sc_hd__clkbuf_2 c69 (.A(net832),
    .X(net49));
 sky130_fd_sc_hd__sdfxtp_1 c690 (.CLK(clknet_leaf_8_clk),
    .D(net685),
    .SCD(net574),
    .SCE(net852),
    .Q(net690));
 sky130_fd_sc_hd__sdfbbn_1 c691 (.CLK_N(clknet_leaf_8_clk),
    .D(net631),
    .RESET_B(net878),
    .SCD(net651),
    .SCE(net688),
    .SET_B(net645),
    .Q(net691));
 sky130_fd_sc_hd__sdfbbp_1 c692 (.CLK(clknet_leaf_8_clk),
    .D(net691),
    .RESET_B(net866),
    .SCD(clknet_1_0__leaf_net535),
    .SCE(net411),
    .SET_B(net864),
    .Q(net692));
 sky130_fd_sc_hd__a21bo_1 c693 (.A1(net532),
    .A2(net13),
    .B1_N(net681),
    .X(net693));
 sky130_fd_sc_hd__clkbuf_1 c694 (.A(net782),
    .X(net694));
 sky130_fd_sc_hd__buf_1 c695 (.A(net782),
    .X(net695));
 sky130_fd_sc_hd__a21bo_1 c696 (.A1(net656),
    .A2(net667),
    .B1_N(net307),
    .X(net696));
 sky130_fd_sc_hd__a21bo_1 c697 (.A1(net424),
    .A2(net694),
    .B1_N(net632),
    .X(net697));
 sky130_fd_sc_hd__sdfxtp_1 c698 (.CLK(clknet_leaf_10_clk),
    .D(net13),
    .SCD(net693),
    .SCE(net191),
    .Q(net698));
 sky130_fd_sc_hd__sdfxtp_1 c699 (.CLK(clknet_leaf_10_clk),
    .D(net584),
    .SCD(net888),
    .SCE(net686),
    .Q(net699));
 sky130_fd_sc_hd__xnor2_1 c70 (.A(net49),
    .B(net834),
    .Y(net50));
 sky130_fd_sc_hd__a21bo_1 c700 (.A1(net679),
    .A2(net672),
    .B1_N(net675),
    .X(net700));
 sky130_fd_sc_hd__xnor2_1 c701 (.A(net836),
    .B(net699),
    .Y(net701));
 sky130_fd_sc_hd__dfbbn_1 c702 (.CLK_N(clknet_leaf_8_clk),
    .D(net654),
    .RESET_B(net666),
    .SET_B(net251),
    .Q(net702));
 sky130_fd_sc_hd__a31o_1 c703 (.A1(net633),
    .A2(net695),
    .A3(net699),
    .B1(net846),
    .X(net703));
 sky130_fd_sc_hd__dfbbn_2 c704 (.CLK_N(clknet_leaf_10_clk),
    .D(net511),
    .RESET_B(net701),
    .SET_B(net664),
    .Q(net705),
    .Q_N(net704));
 sky130_fd_sc_hd__a31o_1 c705 (.A1(net307),
    .A2(net696),
    .A3(net695),
    .B1(net960),
    .X(net706));
 sky130_fd_sc_hd__dfbbp_1 c706 (.CLK(clknet_leaf_14_clk),
    .D(net456),
    .RESET_B(net700),
    .SET_B(net695),
    .Q(net707));
 sky130_fd_sc_hd__a21bo_1 c707 (.A1(net411),
    .A2(net689),
    .B1_N(net696),
    .X(net708));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(net191),
    .A1(net695),
    .A2(net677),
    .A3(net836),
    .S0(net26),
    .S1(net664),
    .X(net709));
 sky130_fd_sc_hd__sedfxbp_1 c709 (.CLK(clknet_leaf_13_clk),
    .D(net561),
    .DE(net708),
    .SCD(net593),
    .SCE(net704),
    .Q(net710));
 sky130_fd_sc_hd__xnor2_4 c71 (.A(net43),
    .B(net798),
    .Y(net51));
 sky130_fd_sc_hd__sdfxbp_1 c710 (.CLK(clknet_leaf_9_clk),
    .D(net650),
    .SCD(net706),
    .SCE(net906),
    .Q(net711));
 sky130_fd_sc_hd__a31o_1 c711 (.A1(net573),
    .A2(net697),
    .A3(net689),
    .B1(net705),
    .X(net712));
 sky130_fd_sc_hd__a21bo_1 c712 (.A1(net707),
    .A2(net710),
    .B1_N(net705),
    .X(net713));
 sky130_fd_sc_hd__sedfxtp_1 c713 (.CLK(clknet_leaf_14_clk),
    .D(net594),
    .DE(net711),
    .SCD(net713),
    .SCE(net664),
    .Q(net714));
 sky130_fd_sc_hd__sedfxtp_1 c714 (.CLK(clknet_leaf_13_clk),
    .D(net397),
    .DE(net705),
    .SCD(net151),
    .SCE(net775),
    .Q(net715));
 sky130_fd_sc_hd__sedfxtp_1 c715 (.CLK(clknet_leaf_14_clk),
    .D(net257),
    .DE(net682),
    .SCD(net895),
    .SCE(net69),
    .Q(net716));
 sky130_fd_sc_hd__a31o_2 c716 (.A1(net11),
    .A2(net676),
    .A3(net475),
    .B1(net593),
    .X(net717));
 sky130_fd_sc_hd__a41o_1 c717 (.A1(net113),
    .A2(net558),
    .A3(net488),
    .A4(net717),
    .B1(net775),
    .X(net718));
 sky130_fd_sc_hd__sdfrbp_1 c718 (.CLK(clknet_leaf_13_clk),
    .D(net69),
    .RESET_B(net562),
    .SCD(net620),
    .SCE(net704),
    .Q(net719));
 sky130_fd_sc_hd__a31o_1 c719 (.A1(net687),
    .A2(net716),
    .A3(net712),
    .B1(net717),
    .X(net720));
 sky130_fd_sc_hd__clkbuf_4 c72 (.A(net755),
    .X(net52));
 sky130_fd_sc_hd__a41o_1 c720 (.A1(net488),
    .A2(net575),
    .A3(net715),
    .A4(net581),
    .B1(net716),
    .X(net721));
 sky130_fd_sc_hd__sdfrbp_1 c721 (.CLK(clknet_leaf_13_clk),
    .D(net516),
    .RESET_B(net858),
    .SCD(net113),
    .SCE(net717),
    .Q(net722));
 sky130_fd_sc_hd__a41o_1 c722 (.A1(net181),
    .A2(net717),
    .A3(net606),
    .A4(net704),
    .B1(net845),
    .X(net723));
 sky130_fd_sc_hd__a41o_1 c723 (.A1(net702),
    .A2(net475),
    .A3(net717),
    .A4(net705),
    .B1(net113),
    .X(net724));
 sky130_fd_sc_hd__sdfrtn_1 c724 (.CLK_N(clknet_leaf_13_clk),
    .D(net721),
    .RESET_B(net847),
    .SCD(net705),
    .SCE(net717),
    .Q(net725));
 sky130_fd_sc_hd__a31o_1 c725 (.A1(net725),
    .A2(net719),
    .A3(net717),
    .B1(net593),
    .X(net726));
 sky130_fd_sc_hd__sdfbbn_1 c726 (.CLK_N(clknet_leaf_13_clk),
    .D(net718),
    .RESET_B(net926),
    .SCD(net682),
    .SCE(net113),
    .SET_B(net939),
    .Q(net727));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net727),
    .A1(net606),
    .A2(net724),
    .A3(net488),
    .S0(net717),
    .S1(net558),
    .X(net728));
 sky130_fd_sc_hd__sdfrtp_1 c728 (.CLK(clknet_leaf_13_clk),
    .D(net893),
    .RESET_B(net664),
    .SCD(net581),
    .SCE(net620),
    .Q(net729));
 sky130_fd_sc_hd__sdfrtp_1 c729 (.CLK(clknet_leaf_13_clk),
    .D(net882),
    .RESET_B(net558),
    .SCD(net726),
    .SCE(net681),
    .Q(net730));
 sky130_fd_sc_hd__buf_1 c73 (.A(net755),
    .X(net53));
 sky130_fd_sc_hd__a31o_1 c730 (.A1(net251),
    .A2(net935),
    .A3(net581),
    .B1(net781),
    .X(net731));
 sky130_fd_sc_hd__sdfrtp_4 c731 (.CLK(clknet_leaf_13_clk),
    .D(net731),
    .RESET_B(net723),
    .SCD(net720),
    .SCE(net676));
 sky130_fd_sc_hd__dfrtp_2 c74 (.CLK(clknet_leaf_31_clk),
    .D(net5),
    .RESET_B(net51),
    .Q(net54));
 sky130_fd_sc_hd__dfrtp_2 c75 (.CLK(clknet_leaf_26_clk),
    .D(net50),
    .RESET_B(net27),
    .Q(net55));
 sky130_fd_sc_hd__dfsbp_1 c76 (.CLK(clknet_leaf_26_clk),
    .D(net916),
    .SET_B(net9),
    .Q(net57),
    .Q_N(net56));
 sky130_fd_sc_hd__xnor2_4 c77 (.A(net49),
    .B(net903),
    .Y(net58));
 sky130_fd_sc_hd__xnor2_1 c78 (.A(net54),
    .B(net11),
    .Y(net59));
 sky130_fd_sc_hd__xnor2_2 c79 (.A(net929),
    .B(net58),
    .Y(net60));
 sky130_fd_sc_hd__xnor2_1 c80 (.A(net58),
    .B(net48),
    .Y(net61));
 sky130_fd_sc_hd__mux4_1 c81 (.A0(net32),
    .A1(net59),
    .A2(net56),
    .A3(net53),
    .S0(net51),
    .S1(net834),
    .X(net62));
 sky130_fd_sc_hd__dfsbp_1 c82 (.CLK(clknet_leaf_25_clk),
    .D(net903),
    .SET_B(net35),
    .Q(net64),
    .Q_N(net63));
 sky130_fd_sc_hd__dfstp_1 c83 (.CLK(clknet_leaf_25_clk),
    .D(net60),
    .SET_B(net61),
    .Q(net65));
 sky130_fd_sc_hd__xnor2_2 c84 (.A(net22),
    .B(net63),
    .Y(net66));
 sky130_fd_sc_hd__clkbuf_4 c85 (.A(net801),
    .X(net67));
 sky130_fd_sc_hd__xnor2_4 c86 (.A(net52),
    .B(net67),
    .Y(net68));
 sky130_fd_sc_hd__xnor2_4 c87 (.A(net28),
    .B(net52),
    .Y(net69));
 sky130_fd_sc_hd__clkbuf_4 c88 (.A(net788),
    .X(net70));
 sky130_fd_sc_hd__xnor2_2 c89 (.A(net955),
    .B(net68),
    .Y(net71));
 sky130_fd_sc_hd__dfstp_1 c90 (.CLK(clknet_leaf_28_clk),
    .D(net787),
    .SET_B(net71),
    .Q(net72));
 sky130_fd_sc_hd__dfstp_1 c91 (.CLK(clknet_leaf_25_clk),
    .D(net35),
    .SET_B(net31),
    .Q(net73));
 sky130_fd_sc_hd__dlrbn_1 c92 (.D(net61),
    .GATE_N(clknet_leaf_25_clk),
    .RESET_B(net801),
    .Q(net75),
    .Q_N(net74));
 sky130_fd_sc_hd__xnor2_2 c93 (.A(net66),
    .B(net70),
    .Y(net76));
 sky130_fd_sc_hd__xnor2_2 c94 (.A(net876),
    .B(net67),
    .Y(net77));
 sky130_fd_sc_hd__sdfrbp_1 c95 (.CLK(clknet_leaf_24_clk),
    .D(net67),
    .RESET_B(net77),
    .SCD(net76),
    .SCE(net834),
    .Q(net79),
    .Q_N(net78));
 sky130_fd_sc_hd__dlrbn_1 c96 (.D(net76),
    .GATE_N(clknet_leaf_25_clk),
    .RESET_B(net873),
    .Q(net81),
    .Q_N(net80));
 sky130_fd_sc_hd__xnor2_1 c97 (.A(net68),
    .B(net72),
    .Y(net82));
 sky130_fd_sc_hd__dlrbp_1 c98 (.D(net72),
    .GATE(clknet_leaf_24_clk),
    .RESET_B(net76),
    .Q(net84),
    .Q_N(net83));
 sky130_fd_sc_hd__xnor2_1 c99 (.A(net77),
    .B(net83),
    .Y(net85));
 sky130_fd_sc_hd__sdfsbp_1 merge732 (.CLK(clknet_leaf_25_clk),
    .D(net0),
    .SCD(net28),
    .SCE(net195),
    .SET_B(net80),
    .Q(net733),
    .Q_N(net732));
 sky130_fd_sc_hd__dlrtn_2 merge733 (.D(net96),
    .GATE_N(clknet_leaf_24_clk),
    .RESET_B(net94),
    .Q(net734));
 sky130_fd_sc_hd__dlrtn_1 merge734 (.D(net253),
    .GATE_N(clknet_leaf_4_clk),
    .RESET_B(net256),
    .Q(net735));
 sky130_fd_sc_hd__dlrtp_1 merge735 (.D(net19),
    .GATE(clknet_leaf_30_clk),
    .RESET_B(clknet_1_1__leaf_net154),
    .Q(net736));
 sky130_fd_sc_hd__dlrtp_1 merge736 (.D(net130),
    .GATE(clknet_leaf_33_clk),
    .RESET_B(net123),
    .Q(net737));
 sky130_fd_sc_hd__sdfsbp_1 merge737 (.CLK(clknet_leaf_17_clk),
    .D(net360),
    .SCD(net604),
    .SCE(net362),
    .SET_B(net490),
    .Q(net739),
    .Q_N(net738));
 sky130_fd_sc_hd__sdfstp_1 merge738 (.CLK(clknet_leaf_17_clk),
    .D(net467),
    .SCD(net405),
    .SCE(net206),
    .SET_B(net360),
    .Q(net740));
 sky130_fd_sc_hd__mux4_1 merge739 (.A0(net677),
    .A1(net692),
    .A2(net26),
    .A3(clknet_1_1__leaf_net535),
    .S0(net683),
    .S1(net532),
    .X(net741));
 sky130_fd_sc_hd__dlrtp_1 merge740 (.D(net9),
    .GATE(clknet_leaf_26_clk),
    .RESET_B(net790),
    .Q(net742));
 sky130_fd_sc_hd__sdfstp_1 merge741 (.CLK(clknet_leaf_12_clk),
    .D(clknet_1_1__leaf_net294),
    .SCD(net516),
    .SCE(net898),
    .SET_B(net582),
    .Q(net743));
 sky130_fd_sc_hd__sdfxbp_1 merge742 (.CLK(clknet_leaf_2_clk),
    .D(net125),
    .SCD(net534),
    .SCE(net151),
    .Q(net745),
    .Q_N(net744));
 sky130_fd_sc_hd__sdfstp_1 merge743 (.CLK(clknet_leaf_12_clk),
    .D(net328),
    .SCD(net950),
    .SCE(net453),
    .SET_B(net961),
    .Q(net746));
 sky130_fd_sc_hd__sdfxtp_1 merge744 (.CLK(clknet_leaf_35_clk),
    .D(clknet_1_1__leaf_net269),
    .SCD(net125),
    .SCE(net419),
    .Q(net747));
 sky130_fd_sc_hd__sedfxbp_1 merge745 (.CLK(clknet_leaf_33_clk),
    .D(net114),
    .DE(net123),
    .SCD(net125),
    .SCE(net124),
    .Q(net749),
    .Q_N(net748));
 sky130_fd_sc_hd__sedfxbp_1 merge746 (.CLK(clknet_leaf_33_clk),
    .D(net8),
    .DE(net119),
    .SCD(clknet_1_0__leaf_net134),
    .SCE(net9),
    .Q(net751),
    .Q_N(net750));
 sky130_fd_sc_hd__mux4_1 merge747 (.A0(net322),
    .A1(net515),
    .A2(net664),
    .A3(net795),
    .S0(net631),
    .S1(net645),
    .X(net752));
 sky130_fd_sc_hd__sedfxtp_1 merge748 (.CLK(clknet_leaf_0_clk),
    .D(net413),
    .DE(net318),
    .SCD(net310),
    .SCE(net799),
    .Q(net753));
 sky130_fd_sc_hd__mux4_1 merge749 (.A0(clknet_1_0__leaf_net372),
    .A1(net823),
    .A2(net236),
    .A3(net795),
    .S0(net414),
    .S1(net776),
    .X(net754));
 sky130_fd_sc_hd__sedfxtp_1 merge750 (.CLK(clknet_leaf_26_clk),
    .D(net42),
    .DE(net51),
    .SCD(net48),
    .SCE(net50),
    .Q(net755));
 sky130_fd_sc_hd__dfxtp_2 s751 (.CLK(clknet_leaf_32_clk),
    .D(net1),
    .Q(net756));
 sky130_fd_sc_hd__dlclkp_1 s752 (.CLK(clknet_leaf_26_clk),
    .GATE(net62),
    .GCLK(net757));
 sky130_fd_sc_hd__dlclkp_2 s753 (.CLK(clknet_leaf_34_clk),
    .GATE(net129),
    .GCLK(net758));
 sky130_fd_sc_hd__dlclkp_4 s754 (.CLK(clknet_leaf_31_clk),
    .GATE(net172),
    .GCLK(net759));
 sky130_fd_sc_hd__dlxbn_1 s755 (.D(net247),
    .GATE_N(clknet_leaf_21_clk),
    .Q(net761),
    .Q_N(net760));
 sky130_fd_sc_hd__dlxbn_1 s756 (.D(net341),
    .GATE_N(clknet_leaf_18_clk),
    .Q(net762));
 sky130_fd_sc_hd__dlxbp_1 s757 (.D(net346),
    .GATE(clknet_leaf_19_clk),
    .Q(net764),
    .Q_N(net763));
 sky130_fd_sc_hd__dlxtn_1 s758 (.D(net364),
    .GATE_N(clknet_leaf_17_clk),
    .Q(net765));
 sky130_fd_sc_hd__dlxtn_1 s759 (.D(net430),
    .GATE_N(clknet_leaf_3_clk),
    .Q(net766));
 sky130_fd_sc_hd__dlxtn_1 s760 (.D(net431),
    .GATE_N(clknet_leaf_3_clk),
    .Q(net767));
 sky130_fd_sc_hd__dlxtp_1 s761 (.D(net446),
    .GATE(clknet_leaf_1_clk),
    .Q(net768));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s762 (.D(net447),
    .SLEEP_B(clknet_leaf_1_clk),
    .Q(net769));
 sky130_fd_sc_hd__dfxbp_1 s763 (.CLK(clknet_leaf_10_clk),
    .D(net452),
    .Q(net771),
    .Q_N(net770));
 sky130_fd_sc_hd__dfxbp_1 s764 (.CLK(clknet_leaf_19_clk),
    .D(net492),
    .Q(net772));
 sky130_fd_sc_hd__dfxtp_1 s765 (.CLK(clknet_leaf_17_clk),
    .D(net494),
    .Q(net773));
 sky130_fd_sc_hd__dfxtp_1 s766 (.CLK(clknet_leaf_13_clk),
    .D(net495),
    .Q(net774));
 sky130_fd_sc_hd__dfxtp_2 s767 (.CLK(clknet_leaf_17_clk),
    .D(net496),
    .Q(net775));
 sky130_fd_sc_hd__dlclkp_1 s768 (.CLK(clknet_leaf_16_clk),
    .GATE(net498),
    .GCLK(net776));
 sky130_fd_sc_hd__dlclkp_2 s769 (.CLK(clknet_leaf_20_clk),
    .GATE(net507),
    .GCLK(net815));
 sky130_fd_sc_hd__dlclkp_4 s770 (.CLK(clknet_leaf_2_clk),
    .GATE(net550),
    .GCLK(net777));
 sky130_fd_sc_hd__dlxbn_1 s771 (.D(net600),
    .GATE_N(clknet_leaf_13_clk),
    .Q(net778));
 sky130_fd_sc_hd__dlxbn_1 s772 (.D(net647),
    .GATE_N(clknet_leaf_7_clk),
    .Q(net779));
 sky130_fd_sc_hd__dlxbp_1 s773 (.D(net709),
    .GATE(clknet_leaf_9_clk),
    .Q(net780));
 sky130_fd_sc_hd__dlxtn_1 s774 (.D(net728),
    .GATE_N(clknet_2_3__leaf_clk),
    .Q(net781));
 sky130_fd_sc_hd__dlxtn_1 s775 (.D(net741),
    .GATE_N(clknet_leaf_9_clk),
    .Q(net782));
 sky130_fd_sc_hd__dlxtn_1 s776 (.D(net752),
    .GATE_N(clknet_leaf_8_clk),
    .Q(net783));
 sky130_fd_sc_hd__dlxtp_1 s777 (.D(net754),
    .GATE(clknet_leaf_16_clk),
    .Q(net784));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(in0),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_8 input2 (.A(in1),
    .X(net786));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(net867),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(in11),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(in12),
    .X(net789));
 sky130_fd_sc_hd__buf_1 input6 (.A(in13),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(in15),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(in16),
    .X(net792));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(in17),
    .X(net793));
 sky130_fd_sc_hd__buf_2 input10 (.A(in18),
    .X(net794));
 sky130_fd_sc_hd__clkbuf_8 input11 (.A(in19),
    .X(net795));
 sky130_fd_sc_hd__buf_4 input12 (.A(in2),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(in20),
    .X(net797));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(in21),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(in22),
    .X(net799));
 sky130_fd_sc_hd__buf_2 input16 (.A(in23),
    .X(net800));
 sky130_fd_sc_hd__buf_4 input17 (.A(in24),
    .X(net801));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(in3),
    .X(net802));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(in4),
    .X(net803));
 sky130_fd_sc_hd__buf_2 input20 (.A(in5),
    .X(net804));
 sky130_fd_sc_hd__buf_4 input21 (.A(in6),
    .X(net805));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(in7),
    .X(net806));
 sky130_fd_sc_hd__buf_2 input23 (.A(in8),
    .X(net807));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(in9),
    .X(net808));
 sky130_fd_sc_hd__buf_2 output25 (.A(net839),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output26 (.A(net810),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output27 (.A(net811),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output28 (.A(net812),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_4 output29 (.A(net813),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output30 (.A(net814),
    .X(out13));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net815),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output32 (.A(net816),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output33 (.A(net817),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output34 (.A(net818),
    .X(out17));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(clknet_1_1__leaf_net819),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output36 (.A(net820),
    .X(out19));
 sky130_fd_sc_hd__clkbuf_4 output37 (.A(net821),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output38 (.A(net822),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output39 (.A(net823),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output40 (.A(net824),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output41 (.A(net825),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output42 (.A(net826),
    .X(out24));
 sky130_fd_sc_hd__clkbuf_1 output43 (.A(clknet_1_1__leaf_net827),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output44 (.A(net828),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output45 (.A(net829),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output46 (.A(net830),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_4 output47 (.A(net831),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output48 (.A(net832),
    .X(out8));
 sky130_fd_sc_hd__clkbuf_1 output49 (.A(net833),
    .X(out9));
 sky130_fd_sc_hd__buf_4 fanout50 (.A(net47),
    .X(net834));
 sky130_fd_sc_hd__buf_4 max_cap51 (.A(net2),
    .X(net835));
 sky130_fd_sc_hd__buf_4 max_cap52 (.A(net122),
    .X(net836));
 sky130_fd_sc_hd__buf_4 max_cap53 (.A(net117),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net759 (.A(net759),
    .X(clknet_0_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net759 (.A(clknet_0_net759),
    .X(clknet_1_0__leaf_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net759 (.A(clknet_0_net759),
    .X(clknet_1_1__leaf_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net176 (.A(net176),
    .X(clknet_0_net176));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net176 (.A(clknet_0_net176),
    .X(clknet_1_0__leaf_net176));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net176 (.A(clknet_0_net176),
    .X(clknet_1_1__leaf_net176));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net174 (.A(net174),
    .X(clknet_0_net174));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net174 (.A(clknet_0_net174),
    .X(clknet_1_0__leaf_net174));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net174 (.A(clknet_0_net174),
    .X(clknet_1_1__leaf_net174));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net758 (.A(net758),
    .X(clknet_0_net758));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net758 (.A(clknet_0_net758),
    .X(clknet_1_0__leaf_net758));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net758 (.A(clknet_0_net758),
    .X(clknet_1_1__leaf_net758));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net400 (.A(net400),
    .X(clknet_0_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net400 (.A(clknet_0_net400),
    .X(clknet_1_0__leaf_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net400 (.A(clknet_0_net400),
    .X(clknet_1_1__leaf_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net401 (.A(net401),
    .X(clknet_0_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net401 (.A(clknet_0_net401),
    .X(clknet_1_0__leaf_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net401 (.A(clknet_0_net401),
    .X(clknet_1_1__leaf_net401));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net421 (.A(net421),
    .X(clknet_0_net421));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net421 (.A(clknet_0_net421),
    .X(clknet_1_0__leaf_net421));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net421 (.A(clknet_0_net421),
    .X(clknet_1_1__leaf_net421));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net398 (.A(net398),
    .X(clknet_0_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_0__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_1__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net269 (.A(net269),
    .X(clknet_0_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net269 (.A(clknet_0_net269),
    .X(clknet_1_0__leaf_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net269 (.A(clknet_0_net269),
    .X(clknet_1_1__leaf_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net757 (.A(net757),
    .X(clknet_0_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net757 (.A(clknet_0_net757),
    .X(clknet_1_0__leaf_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net757 (.A(clknet_0_net757),
    .X(clknet_1_1__leaf_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net250 (.A(net250),
    .X(clknet_0_net250));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net250 (.A(clknet_0_net250),
    .X(clknet_1_0__leaf_net250));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net250 (.A(clknet_0_net250),
    .X(clknet_1_1__leaf_net250));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net827 (.A(net827),
    .X(clknet_0_net827));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net827 (.A(clknet_0_net827),
    .X(clknet_1_0__leaf_net827));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net827 (.A(clknet_0_net827),
    .X(clknet_1_1__leaf_net827));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net205 (.A(net205),
    .X(clknet_0_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net205 (.A(clknet_0_net205),
    .X(clknet_1_0__leaf_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net205 (.A(clknet_0_net205),
    .X(clknet_1_1__leaf_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net103 (.A(net103),
    .X(clknet_0_net103));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net103 (.A(clknet_0_net103),
    .X(clknet_1_0__leaf_net103));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net103 (.A(clknet_0_net103),
    .X(clknet_1_1__leaf_net103));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net108 (.A(net108),
    .X(clknet_0_net108));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net108 (.A(clknet_0_net108),
    .X(clknet_1_0__leaf_net108));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net108 (.A(clknet_0_net108),
    .X(clknet_1_1__leaf_net108));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net274 (.A(net274),
    .X(clknet_0_net274));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net274 (.A(clknet_0_net274),
    .X(clknet_1_0__leaf_net274));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net274 (.A(clknet_0_net274),
    .X(clknet_1_1__leaf_net274));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net293 (.A(net293),
    .X(clknet_0_net293));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net293 (.A(clknet_0_net293),
    .X(clknet_1_0__leaf_net293));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net293 (.A(clknet_0_net293),
    .X(clknet_1_1__leaf_net293));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net280 (.A(net280),
    .X(clknet_0_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net280 (.A(clknet_0_net280),
    .X(clknet_1_0__leaf_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net280 (.A(clknet_0_net280),
    .X(clknet_1_1__leaf_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net294 (.A(net294),
    .X(clknet_0_net294));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net294 (.A(clknet_0_net294),
    .X(clknet_1_0__leaf_net294));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net294 (.A(clknet_0_net294),
    .X(clknet_1_1__leaf_net294));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net264 (.A(net264),
    .X(clknet_0_net264));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net264 (.A(clknet_0_net264),
    .X(clknet_1_0__leaf_net264));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net264 (.A(clknet_0_net264),
    .X(clknet_1_1__leaf_net264));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net303 (.A(net303),
    .X(clknet_0_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net303 (.A(clknet_0_net303),
    .X(clknet_1_0__leaf_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net303 (.A(clknet_0_net303),
    .X(clknet_1_1__leaf_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net443 (.A(net443),
    .X(clknet_0_net443));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net443 (.A(clknet_0_net443),
    .X(clknet_1_0__leaf_net443));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net443 (.A(clknet_0_net443),
    .X(clknet_1_1__leaf_net443));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net451 (.A(net451),
    .X(clknet_0_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net451 (.A(clknet_0_net451),
    .X(clknet_1_0__leaf_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net451 (.A(clknet_0_net451),
    .X(clknet_1_1__leaf_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net448 (.A(net448),
    .X(clknet_0_net448));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net448 (.A(clknet_0_net448),
    .X(clknet_1_0__leaf_net448));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net448 (.A(clknet_0_net448),
    .X(clknet_1_1__leaf_net448));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net435 (.A(net435),
    .X(clknet_0_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net435 (.A(clknet_0_net435),
    .X(clknet_1_0__leaf_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net435 (.A(clknet_0_net435),
    .X(clknet_1_1__leaf_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net272 (.A(net272),
    .X(clknet_0_net272));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net272 (.A(clknet_0_net272),
    .X(clknet_1_0__leaf_net272));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net272 (.A(clknet_0_net272),
    .X(clknet_1_1__leaf_net272));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net262 (.A(net262),
    .X(clknet_0_net262));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net262 (.A(clknet_0_net262),
    .X(clknet_1_0__leaf_net262));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net262 (.A(clknet_0_net262),
    .X(clknet_1_1__leaf_net262));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net292 (.A(net292),
    .X(clknet_0_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net292 (.A(clknet_0_net292),
    .X(clknet_1_0__leaf_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net292 (.A(clknet_0_net292),
    .X(clknet_1_1__leaf_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net267 (.A(net267),
    .X(clknet_0_net267));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net267 (.A(clknet_0_net267),
    .X(clknet_1_0__leaf_net267));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net267 (.A(clknet_0_net267),
    .X(clknet_1_1__leaf_net267));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net521 (.A(net521),
    .X(clknet_0_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net521 (.A(clknet_0_net521),
    .X(clknet_1_0__leaf_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net521 (.A(clknet_0_net521),
    .X(clknet_1_1__leaf_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net268 (.A(net268),
    .X(clknet_0_net268));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net268 (.A(clknet_0_net268),
    .X(clknet_1_0__leaf_net268));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net268 (.A(clknet_0_net268),
    .X(clknet_1_1__leaf_net268));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net265 (.A(net265),
    .X(clknet_0_net265));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net265 (.A(clknet_0_net265),
    .X(clknet_1_0__leaf_net265));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net265 (.A(clknet_0_net265),
    .X(clknet_1_1__leaf_net265));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net287 (.A(net287),
    .X(clknet_0_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net287 (.A(clknet_0_net287),
    .X(clknet_1_0__leaf_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net287 (.A(clknet_0_net287),
    .X(clknet_1_1__leaf_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net139 (.A(net139),
    .X(clknet_0_net139));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net139 (.A(clknet_0_net139),
    .X(clknet_1_0__leaf_net139));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net139 (.A(clknet_0_net139),
    .X(clknet_1_1__leaf_net139));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net143 (.A(net143),
    .X(clknet_0_net143));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net143 (.A(clknet_0_net143),
    .X(clknet_1_0__leaf_net143));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net143 (.A(clknet_0_net143),
    .X(clknet_1_1__leaf_net143));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net187 (.A(net187),
    .X(clknet_0_net187));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net187 (.A(clknet_0_net187),
    .X(clknet_1_0__leaf_net187));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net187 (.A(clknet_0_net187),
    .X(clknet_1_1__leaf_net187));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net204 (.A(net204),
    .X(clknet_0_net204));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net204 (.A(clknet_0_net204),
    .X(clknet_1_0__leaf_net204));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net204 (.A(clknet_0_net204),
    .X(clknet_1_1__leaf_net204));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net202 (.A(net202),
    .X(clknet_0_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net202 (.A(clknet_0_net202),
    .X(clknet_1_0__leaf_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net202 (.A(clknet_0_net202),
    .X(clknet_1_1__leaf_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net147 (.A(net147),
    .X(clknet_0_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net147 (.A(clknet_0_net147),
    .X(clknet_1_0__leaf_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net147 (.A(clknet_0_net147),
    .X(clknet_1_1__leaf_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net142 (.A(net142),
    .X(clknet_0_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net142 (.A(clknet_0_net142),
    .X(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net142 (.A(clknet_0_net142),
    .X(clknet_1_1__leaf_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net535 (.A(net535),
    .X(clknet_0_net535));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net535 (.A(clknet_0_net535),
    .X(clknet_1_0__leaf_net535));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net535 (.A(clknet_0_net535),
    .X(clknet_1_1__leaf_net535));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net279 (.A(net279),
    .X(clknet_0_net279));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net279 (.A(clknet_0_net279),
    .X(clknet_1_0__leaf_net279));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net279 (.A(clknet_0_net279),
    .X(clknet_1_1__leaf_net279));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net148 (.A(net148),
    .X(clknet_0_net148));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net148 (.A(clknet_0_net148),
    .X(clknet_1_0__leaf_net148));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net148 (.A(clknet_0_net148),
    .X(clknet_1_1__leaf_net148));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net146 (.A(net146),
    .X(clknet_0_net146));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net146 (.A(clknet_0_net146),
    .X(clknet_1_0__leaf_net146));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net146 (.A(clknet_0_net146),
    .X(clknet_1_1__leaf_net146));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net134 (.A(net134),
    .X(clknet_0_net134));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net134 (.A(clknet_0_net134),
    .X(clknet_1_0__leaf_net134));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net134 (.A(clknet_0_net134),
    .X(clknet_1_1__leaf_net134));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net154 (.A(net154),
    .X(clknet_0_net154));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net154 (.A(clknet_0_net154),
    .X(clknet_1_0__leaf_net154));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net154 (.A(clknet_0_net154),
    .X(clknet_1_1__leaf_net154));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net112 (.A(net112),
    .X(clknet_0_net112));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net112 (.A(clknet_0_net112),
    .X(clknet_1_0__leaf_net112));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net112 (.A(clknet_0_net112),
    .X(clknet_1_1__leaf_net112));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net372 (.A(net372),
    .X(clknet_0_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_0__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_1__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net819 (.A(net819),
    .X(clknet_0_net819));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net819 (.A(clknet_0_net819),
    .X(clknet_1_0__leaf_net819));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net819 (.A(clknet_0_net819),
    .X(clknet_1_1__leaf_net819));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net234 (.A(net234),
    .X(clknet_0_net234));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net234 (.A(clknet_0_net234),
    .X(clknet_1_0__leaf_net234));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net234 (.A(clknet_0_net234),
    .X(clknet_1_1__leaf_net234));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net239 (.A(net239),
    .X(clknet_0_net239));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net239 (.A(clknet_0_net239),
    .X(clknet_1_0__leaf_net239));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net239 (.A(clknet_0_net239),
    .X(clknet_1_1__leaf_net239));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net233 (.A(net233),
    .X(clknet_0_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net233 (.A(clknet_0_net233),
    .X(clknet_1_0__leaf_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net233 (.A(clknet_0_net233),
    .X(clknet_1_1__leaf_net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net491),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net275),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net309),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net38),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net774),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net778),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net703),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net166),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net178),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net20),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net768),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net771),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net557),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net571),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net529),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net304),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net577),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net581),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net444),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net388),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net157),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net282),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net349),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net770),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net326),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net690),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(in10),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net182),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net420),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net582),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net152),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net235),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net78),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net440),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net153),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net75),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net331),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net680),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net83),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net162),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net261),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net729),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net210),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net426),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net81),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net173),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net305),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net698),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net363),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net576),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net86),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net508),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net722),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net736),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net714),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net772),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net156),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net569),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net322),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net107),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net72),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net348),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net55),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net283),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net463),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net780),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net368),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net248),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net271),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net73),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net522),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net541),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net673),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net553),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net306),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net54),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net155),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net185),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net220),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net34),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net160),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net302),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net566),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net738),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net594),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net593),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(net632),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net41),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net57),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(net590),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net23),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(net402),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(net311),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(net192),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(net730),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(net671),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(net668),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(net591),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(net704),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(net16),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(net674),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(net137),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(net489),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(net652),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(net199),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(net585),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(net635),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(net89),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(net222),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(net428),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(net629),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(net474),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(net352),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(net743),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(net64),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(net628),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(net659),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(net217),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(net316),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(net699),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(net459),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(net330),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(net198),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(net288),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(net739),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(net773),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(net763),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(net768),
    .X(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold30_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge732_D (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c56_RESET_B (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_A3 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c25_Y (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A3 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_SET_B (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_SET_B (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_RESET_B (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_D (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c54_A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_B1_N (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_X (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_SCD (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_SCE (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_SCD (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_B1_N (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A3 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_X (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap53_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_SCD (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_SCD (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_Y (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c642_B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c638_RESET_B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_X (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge746_DE (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_D (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_RESET_B (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_S0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_RESET_B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_D (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_Y (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_D (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_S1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_RESET_B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_X (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap52_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_RESET_B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_RESET_B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_SCE (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_Y (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge745_SCE (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A0 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_X (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge745_SCD (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge744_SCD (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge742_D (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_X (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_D (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_SET_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_X (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_S1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_Y (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_SCD (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_A3 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_SCD (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_B1_N (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_D (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_X (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold105_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_D (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_SCD (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_B (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_Y (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_D (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_SCD (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_RESET_B (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_B1_N (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_Y (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_B (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c54_B1_N (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_X (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A0 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_SCD (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_Q (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge742_SCE (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_SCD (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_GATE (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_RESET_B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_RESET_B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_RESET_B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_X (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold24_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_S1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_Q (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_D (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_SET_B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_SCE (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_X (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_SCE (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_Q_N (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_SCD (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_SCD (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_Q (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_Q (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_SCE (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_SET_B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_Y (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold108_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_Q (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge738_SCE (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_D (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_Y (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_RESET_B (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_SCE (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_SCD (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_DE (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_SCE (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_SCE (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_RESET_B (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_Y (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold121_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_SCD (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A2 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_B1_N (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_Q (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_D (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_X (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c47_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c46_Q (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_SET_B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_SCE (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_SCD (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_X (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_D (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_SET_B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A3 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A3 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_SCD (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_RESET_B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_D (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_Y (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge734_D (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c650_SET_B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c643_D (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_SET_B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_SET_B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_Y (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_RESET_B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_X (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_D (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_B1_N (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_SCD (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_X (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge739_A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c48_Q_N (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_SET_B (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c638_SET_B (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_B (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_GATE (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_Y (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_GATE (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_X (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_RESET_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c51_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c49_Y (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_B1_N (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A3 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_RESET_B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_Y (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold25_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_Q (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_D (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_SCD (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_Q (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_D (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_SCE (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c51_Y (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_SCD (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_Q_N (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_RESET_B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_Q (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_DE (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_B1_N (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_Q (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_B1_N (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_B (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_RESET_B (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_RESET_B (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_X (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_SET_B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c53_X (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_RESET_B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S0 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_B1_N (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_RESET_B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_S0 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_Q (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge748_DE (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_D (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_RESET_B (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_S0 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_RESET_B (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_Y (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A3 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_B1_N (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_Q_N (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_B1_N (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_Q (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold62_A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge747_A0 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A2 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A2 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_Y (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold83_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c61_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c56_Q (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B1_N (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_B1_N (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c58_Y (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_SCD (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_S1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B1_N (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge738_SET_B (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge737_D (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_SCE (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S0 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A3 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_SCD (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_SCD (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_Y (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold23_A (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_Q (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_D (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_RESET_B (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_RESET_B (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_SCD (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_B (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_RESET_B (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_X (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_D (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_B (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_B1_N (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A2 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_B (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_Y (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_B (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_B (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_Q (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c649_D (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_SET_B (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_SCE (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_Y (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge738_SCD (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_Q_N (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_Q (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_RESET_B (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_B (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_Q_N (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A2 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_Q (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_SCE (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_SCE (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_SCD (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A3 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A3 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_B1_N (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_Y (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge749_S0 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_D (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_SET_B (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A3 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_S0 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_SCD (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_SET_B (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_Y (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_B (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A2 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_Q (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold113_A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_RESET_B (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_B1 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_B1_N (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_Q (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A3 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_X (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_D (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_SCD (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_Q (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_D (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_B1_N (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_Y (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A3 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_SCD (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A3 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_Y (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4_A (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_B1_N (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_B1_N (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A2 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_Q (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_D (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c39_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c30_X (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge750_DE (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_S0 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_RESET_B (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_Y (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_RESET_B (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_D (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_RESET_B (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A1 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_B1 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_SET_B (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_X (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_D (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_c657_SCE (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_RESET_B (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_B (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_B (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_X (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge747_A1 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_B1_N (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A4 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_D (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_RESET_B (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_B (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_X (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge741_SCD (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_D (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_SCD (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_RESET_B (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_S1 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_Y (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_SCE (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_SCE (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_B (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_Q (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge739_S1 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A1 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A3 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A3 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A2 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_X (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold79_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_Q (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_B1_N (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_S1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_Q (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold75_A (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_B (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_Q (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A0 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_SCE (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A3 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_X (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_Q (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_RESET_B (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A2 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_B1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_Y (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_GCLK (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold33_A (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge741_SET_B (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_D (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_SCD (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_X (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_SET_B (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_D (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_Y (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge747_S0 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_D (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_D (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c641_SET_B (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c640_Y (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold90_A (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_B1_N (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_B1_N (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c641_Q_N (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A1 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_B1_N (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c649_SCD (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c641_Q (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge747_S1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_SET_B (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_D (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_RESET_B (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_RESET_B (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_SET_B (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c653_RESET_B (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c652_Y (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge747_A2 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_RESET_B (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_SCE (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_SET_B (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_SCD (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_RESET_B (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_SCE (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_Y (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_SCE (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_Q (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_SCD (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_DE (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_SCE (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_Q (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_Y (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_D (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_SCE (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_SET_B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_SCE (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_RESET_B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_D (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_SCE (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_Q (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_s751_Q (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_B (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_SET_B (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_B (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_s767_Q (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_B1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_SCE (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_SET_B (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_B1_N (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_SET_B (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge746_SCE (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge740_D (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_SET_B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_Y (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_D (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_D (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_D (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_X (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_A2 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_D (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_B1_N (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_D (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_B (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_RESET_B (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A2 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_B1_N (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c53_A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c35_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_B (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_B (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c28_A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge749_A3 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge747_A3 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_B1_N (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_B (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_B (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c54_A2 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge748_SCE (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_RESET_B (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A3 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_A0 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_B1_N (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_RESET_B (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c58_B (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c27_A (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A0 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c58_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_SET_B (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_D (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_SCE (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_output25_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_B1_N (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A3 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_B1_N (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_X (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_output29_A (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_RESET_B (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_SCD (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_SCE (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_X (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_output32_A (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A3 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_B1_N (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B1_N (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A2 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_SET_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_RESET_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A2 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_Q (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_output39_A (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge749_A1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A3 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A3 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_SET_B (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_Q (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_SCE (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_Y (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_output48_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_SET_B (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c48_Q (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_B1_N (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_D (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_X (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_SCD (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_SCE (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_SCE (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_B1_N (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_B1_N (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_S1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_B (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_B1_N (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A3 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap51_X (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_B (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap52_X (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_S1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A3 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge741_CLK (.DIODE(clknet_leaf_12_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_CLK (.DIODE(clknet_leaf_12_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_CLK (.DIODE(clknet_leaf_12_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_GATE_N (.DIODE(clknet_leaf_12_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_CLK (.DIODE(clknet_leaf_12_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_CLK_N (.DIODE(clknet_leaf_12_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge743_CLK (.DIODE(clknet_leaf_12_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_GATE_N (.DIODE(clknet_leaf_12_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_CLK (.DIODE(clknet_leaf_12_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_CLK (.DIODE(clknet_leaf_12_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_CLK (.DIODE(clknet_leaf_12_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_CLK (.DIODE(clknet_leaf_12_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_CLK (.DIODE(clknet_leaf_12_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_X (.DIODE(clknet_leaf_12_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_CLK_N (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_GATE_N (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_CLK (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_CLK (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_GATE (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_CLK_N (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_GATE (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_CLK (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_GATE (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_CLK (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_CLK_N (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_GATE_N (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_GATE (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_X (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_X (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_X (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_X (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s774_GATE_N (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_X (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_RESET_B (.DIODE(clknet_1_0__leaf_net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_RESET_B (.DIODE(clknet_1_0__leaf_net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_RESET_B (.DIODE(clknet_1_0__leaf_net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net294_X (.DIODE(clknet_1_0__leaf_net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_SCE (.DIODE(clknet_1_1__leaf_net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_SET_B (.DIODE(clknet_1_1__leaf_net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_SET_B (.DIODE(clknet_1_1__leaf_net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge741_D (.DIODE(clknet_1_1__leaf_net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net294_X (.DIODE(clknet_1_1__leaf_net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_SCE (.DIODE(clknet_1_1__leaf_net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_RESET_B (.DIODE(clknet_1_1__leaf_net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_D (.DIODE(clknet_1_1__leaf_net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net187_X (.DIODE(clknet_1_1__leaf_net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_RESET_B (.DIODE(clknet_1_0__leaf_net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_SET_B (.DIODE(clknet_1_0__leaf_net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S1 (.DIODE(clknet_1_0__leaf_net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_SCE (.DIODE(clknet_1_0__leaf_net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_SCE (.DIODE(clknet_1_0__leaf_net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S1 (.DIODE(clknet_1_0__leaf_net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net202_X (.DIODE(clknet_1_0__leaf_net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_RESET_B (.DIODE(clknet_1_1__leaf_net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_SCE (.DIODE(clknet_1_1__leaf_net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_D (.DIODE(clknet_1_1__leaf_net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net202_X (.DIODE(clknet_1_1__leaf_net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_A (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold23_X (.DIODE(net860));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net237),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net809),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net809),
    .X(net840));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
