module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in3,
    in4,
    in5,
    in6,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out3,
    out4,
    out5,
    out6,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in3;
 input in4;
 input in5;
 input in6;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out3;
 output out4;
 output out5;
 output out6;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net738;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net924;
 wire clknet_1_0__leaf_net924;
 wire clknet_1_1__leaf_net924;
 wire clknet_0_net415;
 wire clknet_1_0__leaf_net415;
 wire clknet_1_1__leaf_net415;
 wire clknet_0_net555;
 wire clknet_1_0__leaf_net555;
 wire clknet_1_1__leaf_net555;
 wire clknet_0_net883;
 wire clknet_1_0__leaf_net883;
 wire clknet_1_1__leaf_net883;
 wire clknet_0_net589;
 wire clknet_1_0__leaf_net589;
 wire clknet_1_1__leaf_net589;
 wire clknet_0_net587;
 wire clknet_1_0__leaf_net587;
 wire clknet_1_1__leaf_net587;
 wire clknet_0_net584;
 wire clknet_1_0__leaf_net584;
 wire clknet_1_1__leaf_net584;
 wire clknet_0_net961;
 wire clknet_1_0__leaf_net961;
 wire clknet_1_1__leaf_net961;
 wire clknet_0_net583;
 wire clknet_1_0__leaf_net583;
 wire clknet_1_1__leaf_net583;
 wire clknet_0_net982;
 wire clknet_1_0__leaf_net982;
 wire clknet_1_1__leaf_net982;
 wire clknet_0_net273;
 wire clknet_1_0__leaf_net273;
 wire clknet_1_1__leaf_net273;
 wire clknet_0_net281;
 wire clknet_1_0__leaf_net281;
 wire clknet_1_1__leaf_net281;
 wire clknet_0_net411;
 wire clknet_1_0__leaf_net411;
 wire clknet_1_1__leaf_net411;
 wire clknet_0_net553;
 wire clknet_1_0__leaf_net553;
 wire clknet_1_1__leaf_net553;
 wire clknet_0_net274;
 wire clknet_1_0__leaf_net274;
 wire clknet_1_1__leaf_net274;
 wire clknet_0_net922;
 wire clknet_1_0__leaf_net922;
 wire clknet_1_1__leaf_net922;
 wire clknet_0_net327;
 wire clknet_1_0__leaf_net327;
 wire clknet_1_1__leaf_net327;
 wire clknet_0_net491;
 wire clknet_1_0__leaf_net491;
 wire clknet_1_1__leaf_net491;
 wire clknet_0_net497;
 wire clknet_1_0__leaf_net497;
 wire clknet_1_1__leaf_net497;
 wire clknet_0_net485;
 wire clknet_1_0__leaf_net485;
 wire clknet_1_1__leaf_net485;
 wire clknet_0_net453;
 wire clknet_1_0__leaf_net453;
 wire clknet_1_1__leaf_net453;
 wire clknet_0_net969;
 wire clknet_1_0__leaf_net969;
 wire clknet_1_1__leaf_net969;
 wire clknet_0_net280;
 wire clknet_1_0__leaf_net280;
 wire clknet_1_1__leaf_net280;
 wire clknet_0_net291;
 wire clknet_1_0__leaf_net291;
 wire clknet_1_1__leaf_net291;
 wire clknet_0_net314;
 wire clknet_1_0__leaf_net314;
 wire clknet_1_1__leaf_net314;
 wire clknet_0_net882;
 wire clknet_1_0__leaf_net882;
 wire clknet_1_1__leaf_net882;
 wire clknet_0_net328;
 wire clknet_1_0__leaf_net328;
 wire clknet_1_1__leaf_net328;
 wire clknet_0_net473;
 wire clknet_1_0__leaf_net473;
 wire clknet_1_1__leaf_net473;
 wire clknet_0_net456;
 wire clknet_1_0__leaf_net456;
 wire clknet_1_1__leaf_net456;
 wire clknet_0_net923;
 wire clknet_1_0__leaf_net923;
 wire clknet_1_1__leaf_net923;
 wire clknet_0_net307;
 wire clknet_1_0__leaf_net307;
 wire clknet_1_1__leaf_net307;
 wire clknet_0_net451;
 wire clknet_1_0__leaf_net451;
 wire clknet_1_1__leaf_net451;
 wire clknet_0_net450;
 wire clknet_1_0__leaf_net450;
 wire clknet_1_1__leaf_net450;
 wire clknet_0_net963;
 wire clknet_1_0__leaf_net963;
 wire clknet_1_1__leaf_net963;
 wire clknet_0_net460;
 wire clknet_1_0__leaf_net460;
 wire clknet_1_1__leaf_net460;
 wire clknet_0_net441;
 wire clknet_1_0__leaf_net441;
 wire clknet_1_1__leaf_net441;
 wire clknet_0_net698;
 wire clknet_1_0__leaf_net698;
 wire clknet_1_1__leaf_net698;
 wire clknet_0_net904;
 wire clknet_1_0__leaf_net904;
 wire clknet_1_1__leaf_net904;
 wire clknet_0_net708;
 wire clknet_1_0__leaf_net708;
 wire clknet_1_1__leaf_net708;
 wire clknet_0_net316;
 wire clknet_1_0__leaf_net316;
 wire clknet_1_1__leaf_net316;
 wire clknet_0_net295;
 wire clknet_1_0__leaf_net295;
 wire clknet_1_1__leaf_net295;
 wire clknet_0_net863;
 wire clknet_1_0__leaf_net863;
 wire clknet_1_1__leaf_net863;
 wire clknet_0_net862;
 wire clknet_1_0__leaf_net862;
 wire clknet_1_1__leaf_net862;
 wire clknet_0_net843;
 wire clknet_1_0__leaf_net843;
 wire clknet_1_1__leaf_net843;
 wire clknet_0_net310;
 wire clknet_1_0__leaf_net310;
 wire clknet_1_1__leaf_net310;
 wire clknet_0_net197;
 wire clknet_1_0__leaf_net197;
 wire clknet_1_1__leaf_net197;
 wire clknet_0_net217;
 wire clknet_1_0__leaf_net217;
 wire clknet_1_1__leaf_net217;
 wire clknet_0_net348;
 wire clknet_1_0__leaf_net348;
 wire clknet_1_1__leaf_net348;
 wire clknet_0_net218;
 wire clknet_1_0__leaf_net218;
 wire clknet_1_1__leaf_net218;
 wire clknet_0_net212;
 wire clknet_1_0__leaf_net212;
 wire clknet_1_1__leaf_net212;
 wire clknet_0_net962;
 wire clknet_1_0__leaf_net962;
 wire clknet_1_1__leaf_net962;
 wire clknet_0_net345;
 wire clknet_1_0__leaf_net345;
 wire clknet_1_1__leaf_net345;
 wire clknet_0_net842;
 wire clknet_1_0__leaf_net842;
 wire clknet_1_1__leaf_net842;
 wire clknet_0_net965;
 wire clknet_1_0__leaf_net965;
 wire clknet_1_1__leaf_net965;
 wire clknet_0_net841;
 wire clknet_1_0__leaf_net841;
 wire clknet_1_1__leaf_net841;
 wire clknet_0_net192;
 wire clknet_1_0__leaf_net192;
 wire clknet_1_1__leaf_net192;
 wire clknet_0_net815;
 wire clknet_1_0__leaf_net815;
 wire clknet_1_1__leaf_net815;
 wire clknet_0_net202;
 wire clknet_1_0__leaf_net202;
 wire clknet_1_1__leaf_net202;
 wire clknet_0_net203;
 wire clknet_1_0__leaf_net203;
 wire clknet_1_1__leaf_net203;
 wire clknet_0_net971;
 wire clknet_1_0__leaf_net971;
 wire clknet_1_1__leaf_net971;
 wire clknet_0_net172;
 wire clknet_1_0__leaf_net172;
 wire clknet_1_1__leaf_net172;
 wire clknet_0_net294;
 wire clknet_1_0__leaf_net294;
 wire clknet_1_1__leaf_net294;
 wire clknet_0_net427;
 wire clknet_1_0__leaf_net427;
 wire clknet_1_1__leaf_net427;
 wire clknet_0_net315;
 wire clknet_1_0__leaf_net315;
 wire clknet_1_1__leaf_net315;
 wire clknet_0_net977;
 wire clknet_1_0__leaf_net977;
 wire clknet_1_1__leaf_net977;
 wire clknet_0_net814;
 wire clknet_1_0__leaf_net814;
 wire clknet_1_1__leaf_net814;
 wire clknet_0_net269;
 wire clknet_1_0__leaf_net269;
 wire clknet_1_1__leaf_net269;
 wire clknet_0_net537;
 wire clknet_1_0__leaf_net537;
 wire clknet_1_1__leaf_net537;
 wire clknet_0_net263;
 wire clknet_1_0__leaf_net263;
 wire clknet_1_1__leaf_net263;
 wire clknet_0_net813;
 wire clknet_1_0__leaf_net813;
 wire clknet_1_1__leaf_net813;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;

 sky130_fd_sc_hd__clkbuf_2 c100 (.A(net782),
    .X(net76));
 sky130_fd_sc_hd__and2_1 c101 (.A(net45),
    .B(net75),
    .X(net77));
 sky130_fd_sc_hd__and2_1 c102 (.A(net72),
    .B(net65),
    .X(net78));
 sky130_fd_sc_hd__and2_0 c103 (.A(net7),
    .B(net75),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 c104 (.A(net1025),
    .X(net80));
 sky130_fd_sc_hd__and2_1 c105 (.A(net80),
    .B(net32),
    .X(net81));
 sky130_fd_sc_hd__sdfbbn_1 c106 (.CLK_N(clknet_4_13_0_clk),
    .D(net44),
    .RESET_B(net79),
    .SCD(net81),
    .SCE(net75),
    .SET_B(net996),
    .Q(net83),
    .Q_N(net82));
 sky130_fd_sc_hd__buf_2 c107 (.A(net781),
    .X(net84));
 sky130_fd_sc_hd__mux4_1 c108 (.A0(net79),
    .A1(net56),
    .A2(net83),
    .A3(net81),
    .S0(net84),
    .S1(net75),
    .X(net85));
 sky130_fd_sc_hd__mux4_1 c109 (.A0(net84),
    .A1(net83),
    .A2(net81),
    .A3(net65),
    .S0(net996),
    .S1(net782),
    .X(net86));
 sky130_fd_sc_hd__and2_1 c110 (.A(net54),
    .B(net837),
    .X(net87));
 sky130_fd_sc_hd__and2_1 c111 (.A(net98),
    .B(net105),
    .X(net88));
 sky130_fd_sc_hd__and2_1 c112 (.A(net27),
    .B(net106),
    .X(net89));
 sky130_fd_sc_hd__mux4_1 c113 (.A0(net104),
    .A1(net89),
    .A2(net87),
    .A3(net65),
    .S0(net71),
    .S1(net70),
    .X(net90));
 sky130_fd_sc_hd__and2_1 c114 (.A(net108),
    .B(net88),
    .X(net91));
 sky130_fd_sc_hd__mux4_1 c115 (.A0(net74),
    .A1(net90),
    .A2(net87),
    .A3(net88),
    .S0(net89),
    .S1(net70),
    .X(net92));
 sky130_fd_sc_hd__and2_0 c116 (.A(net107),
    .B(net91),
    .X(net93));
 sky130_fd_sc_hd__and2_0 c117 (.A(net54),
    .B(net71),
    .X(net94));
 sky130_fd_sc_hd__and2_0 c118 (.A(net75),
    .B(net27),
    .X(net95));
 sky130_fd_sc_hd__and2_0 c119 (.A(net95),
    .B(net27),
    .X(net96));
 sky130_fd_sc_hd__and2_1 c120 (.A(net15),
    .B(net70),
    .X(net97));
 sky130_fd_sc_hd__and2_0 c121 (.A(net97),
    .B(net94),
    .X(net98));
 sky130_fd_sc_hd__and2_1 c122 (.A(net952),
    .B(net27),
    .X(net99));
 sky130_fd_sc_hd__and2_0 c123 (.A(net94),
    .B(net75),
    .X(net100));
 sky130_fd_sc_hd__buf_2 c124 (.A(net807),
    .X(net101));
 sky130_fd_sc_hd__and2_0 c125 (.A(net8),
    .B(net66),
    .X(net102));
 sky130_fd_sc_hd__and2_0 c126 (.A(net99),
    .B(net101),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 c127 (.A(net807),
    .X(net104));
 sky130_fd_sc_hd__or4bb_1 c128 (.A(net103),
    .B(net97),
    .C_N(net101),
    .D_N(net99),
    .X(net105));
 sky130_fd_sc_hd__and2_1 c129 (.A(net96),
    .B(net101),
    .X(net106));
 sky130_fd_sc_hd__and2_0 c130 (.A(net100),
    .B(net105),
    .X(net107));
 sky130_fd_sc_hd__and2_0 c131 (.A(net101),
    .B(net97),
    .X(net108));
 sky130_fd_sc_hd__and2_1 c132 (.A(net944),
    .B(net940),
    .X(net109));
 sky130_fd_sc_hd__and2_1 c133 (.A(net947),
    .B(net109),
    .X(net110));
 sky130_fd_sc_hd__and3_4 c134 (.A(net109),
    .B(net957),
    .C(net945),
    .X(net111));
 sky130_fd_sc_hd__and2_2 c135 (.A(net938),
    .B(net109),
    .X(net112));
 sky130_fd_sc_hd__and2_1 c136 (.A(net112),
    .B(net957),
    .X(net113));
 sky130_fd_sc_hd__and2_1 c137 (.A(net940),
    .B(net109),
    .X(net114));
 sky130_fd_sc_hd__and2_2 c138 (.A(net113),
    .B(net111),
    .X(net115));
 sky130_fd_sc_hd__and2_2 c139 (.A(net738),
    .B(net997),
    .X(net116));
 sky130_fd_sc_hd__and2_1 c140 (.A(net114),
    .B(net947),
    .X(net117));
 sky130_fd_sc_hd__and2_1 c141 (.A(net738),
    .B(net113),
    .X(net118));
 sky130_fd_sc_hd__and2_2 c142 (.A(net940),
    .B(net109),
    .X(net119));
 sky130_fd_sc_hd__and2_1 c143 (.A(net117),
    .B(net119),
    .X(net120));
 sky130_fd_sc_hd__and3_1 c144 (.A(net120),
    .B(net118),
    .C(net117),
    .X(net121));
 sky130_fd_sc_hd__and3_1 c145 (.A(net997),
    .B(net121),
    .C(net118),
    .X(net122));
 sky130_fd_sc_hd__and2_2 c146 (.A(net122),
    .B(net997),
    .X(net123));
 sky130_fd_sc_hd__and2_2 c147 (.A(net110),
    .B(net122),
    .X(net124));
 sky130_fd_sc_hd__and3_4 c148 (.A(net124),
    .B(net113),
    .C(net114),
    .X(net979));
 sky130_fd_sc_hd__and2_4 c149 (.A(net121),
    .B(net114),
    .X(net125));
 sky130_fd_sc_hd__and3_1 c150 (.A(net125),
    .B(net112),
    .C(net123),
    .X(net126));
 sky130_fd_sc_hd__or4bb_2 c151 (.A(net126),
    .B(net125),
    .C_N(net123),
    .D_N(net114),
    .X(net127));
 sky130_fd_sc_hd__mux4_1 c152 (.A0(net127),
    .A1(net111),
    .A2(net110),
    .A3(net118),
    .S0(net121),
    .S1(net997),
    .X(net128));
 sky130_fd_sc_hd__and3_1 c153 (.A(net118),
    .B(net128),
    .C(net127),
    .X(net129));
 sky130_fd_sc_hd__and2_1 c154 (.A(net128),
    .B(net129),
    .X(net130));
 sky130_fd_sc_hd__and2_1 c155 (.A(net128),
    .B(net125),
    .X(net131));
 sky130_fd_sc_hd__and2_1 c156 (.A(net956),
    .B(net131),
    .X(net132));
 sky130_fd_sc_hd__and2_1 c157 (.A(net17),
    .B(net6),
    .X(net133));
 sky130_fd_sc_hd__and2_4 c158 (.A(net951),
    .B(net17),
    .X(net134));
 sky130_fd_sc_hd__and2_4 c159 (.A(net13),
    .B(net979),
    .X(net135));
 sky130_fd_sc_hd__or4bb_1 c160 (.A(net958),
    .B(net133),
    .C_N(net128),
    .D_N(net109),
    .X(net136));
 sky130_fd_sc_hd__and2_1 c161 (.A(net953),
    .B(net129),
    .X(net137));
 sky130_fd_sc_hd__and2_0 c162 (.A(net17),
    .B(net18),
    .X(net138));
 sky130_fd_sc_hd__and2_1 c163 (.A(net138),
    .B(net136),
    .X(net139));
 sky130_fd_sc_hd__and2_0 c164 (.A(net133),
    .B(net138),
    .X(net140));
 sky130_fd_sc_hd__and2_1 c165 (.A(net140),
    .B(net135),
    .X(net141));
 sky130_fd_sc_hd__and2_1 c166 (.A(net137),
    .B(net140),
    .X(net142));
 sky130_fd_sc_hd__and2_2 c167 (.A(net141),
    .B(net132),
    .X(net143));
 sky130_fd_sc_hd__or4bb_1 c168 (.A(net113),
    .B(net141),
    .C_N(net143),
    .D_N(net142),
    .X(net144));
 sky130_fd_sc_hd__sdfrbp_2 c169 (.CLK(clknet_4_5_0_clk),
    .D(net142),
    .RESET_B(net143),
    .SCD(net135),
    .SCE(clknet_1_0__leaf_net815),
    .Q(net146),
    .Q_N(net145));
 sky130_fd_sc_hd__or4bb_1 c170 (.A(net109),
    .B(net131),
    .C_N(net146),
    .D_N(net139),
    .X(net147));
 sky130_fd_sc_hd__mux4_1 c171 (.A0(net143),
    .A1(net140),
    .A2(net147),
    .A3(net146),
    .S0(net135),
    .S1(net18),
    .X(net148));
 sky130_fd_sc_hd__mux4_1 c172 (.A0(net137),
    .A1(net941),
    .A2(net146),
    .A3(net142),
    .S0(net957),
    .S1(clknet_1_0__leaf_net815),
    .X(net977));
 sky130_fd_sc_hd__mux4_1 c173 (.A0(net6),
    .A1(net147),
    .A2(net137),
    .A3(clknet_1_0__leaf_net977),
    .S0(net143),
    .S1(net145),
    .X(net149));
 sky130_fd_sc_hd__sdfrbp_2 c174 (.CLK(clknet_4_5_0_clk),
    .D(net138),
    .RESET_B(net124),
    .SCD(net143),
    .SCE(net833),
    .Q(net151),
    .Q_N(net150));
 sky130_fd_sc_hd__mux4_1 c175 (.A0(net147),
    .A1(net151),
    .A2(net142),
    .A3(net17),
    .S0(net143),
    .S1(net833),
    .X(net152));
 sky130_fd_sc_hd__and2_1 c176 (.A(net945),
    .B(net135),
    .X(net153));
 sky130_fd_sc_hd__and2_2 c177 (.A(net7),
    .B(net833),
    .X(net154));
 sky130_fd_sc_hd__and2_0 c178 (.A(net29),
    .B(net997),
    .X(net155));
 sky130_fd_sc_hd__and2_2 c179 (.A(net16),
    .B(net142),
    .X(net156));
 sky130_fd_sc_hd__and2_0 c180 (.A(net10),
    .B(net125),
    .X(net157));
 sky130_fd_sc_hd__and2_1 c181 (.A(net130),
    .B(net33),
    .X(net158));
 sky130_fd_sc_hd__buf_1 c182 (.A(net731),
    .X(net159));
 sky130_fd_sc_hd__a2111o_1 c183 (.A1(net130),
    .A2(net156),
    .B1(net159),
    .C1(net124),
    .D1(net134),
    .X(net160));
 sky130_fd_sc_hd__sdfrtn_1 c184 (.CLK_N(clknet_4_5_0_clk),
    .D(net153),
    .RESET_B(net24),
    .SCD(net21),
    .SCE(clknet_1_0__leaf_net977),
    .Q(net161));
 sky130_fd_sc_hd__buf_1 c185 (.A(net730),
    .X(net162));
 sky130_fd_sc_hd__and3_2 c186 (.A(net945),
    .B(net6),
    .C(net1037),
    .X(net163));
 sky130_fd_sc_hd__and2_1 c187 (.A(net956),
    .B(net158),
    .X(net164));
 sky130_fd_sc_hd__and2_0 c188 (.A(net154),
    .B(net29),
    .X(net165));
 sky130_fd_sc_hd__and2_0 c189 (.A(net13),
    .B(net154),
    .X(net166));
 sky130_fd_sc_hd__a2111o_1 c190 (.A1(net958),
    .A2(net161),
    .B1(net154),
    .C1(net995),
    .D1(net164),
    .X(net167));
 sky130_fd_sc_hd__a2111o_1 c191 (.A1(net158),
    .A2(net166),
    .B1(net1027),
    .C1(net26),
    .D1(net33),
    .X(net168));
 sky130_fd_sc_hd__sdfrtp_4 c192 (.CLK(clknet_4_5_0_clk),
    .D(net164),
    .RESET_B(net168),
    .SCD(net167),
    .SCE(net145),
    .Q(net981));
 sky130_fd_sc_hd__or4bb_2 c193 (.A(net0),
    .B(net158),
    .C_N(net164),
    .D_N(net24),
    .X(net169));
 sky130_fd_sc_hd__and2_1 c194 (.A(net161),
    .B(net945),
    .X(net170));
 sky130_fd_sc_hd__mux4_1 c195 (.A0(net167),
    .A1(net1006),
    .A2(net164),
    .A3(net169),
    .S0(net168),
    .S1(net1053),
    .X(net171));
 sky130_fd_sc_hd__mux4_1 c196 (.A0(net132),
    .A1(net157),
    .A2(net29),
    .A3(net7),
    .S0(net995),
    .S1(clknet_1_0__leaf_net815),
    .X(net172));
 sky130_fd_sc_hd__mux4_1 c197 (.A0(net142),
    .A1(net1006),
    .A2(net139),
    .A3(net130),
    .S0(net39),
    .S1(net1016),
    .X(net173));
 sky130_fd_sc_hd__and2_1 c198 (.A(net134),
    .B(net155),
    .X(net975));
 sky130_fd_sc_hd__and3_1 c199 (.A(net957),
    .B(net941),
    .C(net953),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 c200 (.A(net914),
    .X(net175));
 sky130_fd_sc_hd__and3_1 c201 (.A(net57),
    .B(net145),
    .C(net788),
    .X(net176));
 sky130_fd_sc_hd__dlymetal6s2s_1 c202 (.A(net914),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 c203 (.A(net1043),
    .X(net178));
 sky130_fd_sc_hd__a2111o_1 c204 (.A1(net177),
    .A2(net56),
    .B1(net51),
    .C1(net986),
    .D1(net1042),
    .X(net179));
 sky130_fd_sc_hd__sdfrtp_1 c205 (.CLK(clknet_4_7_0_clk),
    .D(net116),
    .RESET_B(net49),
    .SCD(net176),
    .SCE(net986),
    .Q(net180));
 sky130_fd_sc_hd__buf_1 c206 (.A(net804),
    .X(net181));
 sky130_fd_sc_hd__sdfbbp_1 c207 (.CLK(clknet_4_13_0_clk),
    .D(net178),
    .RESET_B(net181),
    .SCD(net176),
    .SCE(net986),
    .SET_B(net1017),
    .Q(net183),
    .Q_N(net182));
 sky130_fd_sc_hd__or4bb_1 c208 (.A(net49),
    .B(net57),
    .C_N(net175),
    .D_N(net182),
    .X(net184));
 sky130_fd_sc_hd__a2111o_1 c209 (.A1(net26),
    .A2(net21),
    .B1(net177),
    .C1(net182),
    .D1(net57),
    .X(net185));
 sky130_fd_sc_hd__sdfbbn_1 c210 (.CLK_N(clknet_4_12_0_clk),
    .D(net176),
    .RESET_B(net163),
    .SCD(net180),
    .SCE(net984),
    .SET_B(net937),
    .Q(net187),
    .Q_N(net186));
 sky130_fd_sc_hd__or4bb_1 c211 (.A(net168),
    .B(net177),
    .C_N(net176),
    .D_N(net984),
    .X(net188));
 sky130_fd_sc_hd__mux4_1 c212 (.A0(net174),
    .A1(net184),
    .A2(net26),
    .A3(net984),
    .S0(net176),
    .S1(net181),
    .X(net189));
 sky130_fd_sc_hd__sdfbbn_1 c213 (.CLK_N(clknet_4_13_0_clk),
    .D(net181),
    .RESET_B(net984),
    .SCD(net942),
    .SCE(net36),
    .SET_B(clknet_1_1__leaf_net841),
    .Q(net191),
    .Q_N(net190));
 sky130_fd_sc_hd__mux4_1 c214 (.A0(net174),
    .A1(net178),
    .A2(net57),
    .A3(clknet_1_1__leaf_net813),
    .S0(net840),
    .S1(clknet_1_1__leaf_net841),
    .X(net192));
 sky130_fd_sc_hd__sdfbbp_1 c215 (.CLK(clknet_4_12_0_clk),
    .D(net984),
    .RESET_B(net180),
    .SCD(net190),
    .SCE(clknet_1_0__leaf_net813),
    .SET_B(clknet_1_1__leaf_net841),
    .Q(net194),
    .Q_N(net193));
 sky130_fd_sc_hd__mux4_1 c216 (.A0(net41),
    .A1(net193),
    .A2(net984),
    .A3(net36),
    .S0(net174),
    .S1(clknet_1_0__leaf_net813),
    .X(net195));
 sky130_fd_sc_hd__a2111o_1 c217 (.A1(net132),
    .A2(net183),
    .B1(net49),
    .C1(net986),
    .D1(clknet_1_0__leaf_net842),
    .X(net965));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(net194),
    .A1(net942),
    .A2(clknet_1_1__leaf_net965),
    .A3(net10),
    .S0(net984),
    .S1(clknet_1_1__leaf_net842),
    .X(net196));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net180),
    .A1(net194),
    .A2(net134),
    .A3(clknet_1_1__leaf_net841),
    .S0(clknet_1_1__leaf_net842),
    .S1(clknet_1_1__leaf_net843),
    .X(net197));
 sky130_fd_sc_hd__and2_1 c220 (.A(net155),
    .B(net177),
    .X(net198));
 sky130_fd_sc_hd__or4bb_1 c221 (.A(net10),
    .B(net78),
    .C_N(net76),
    .D_N(net838),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_1 c222 (.A(net808),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_1 c223 (.A(net808),
    .X(net201));
 sky130_fd_sc_hd__and2_0 c224 (.A(clknet_1_1__leaf_net815),
    .B(net839),
    .X(net202));
 sky130_fd_sc_hd__and3_1 c225 (.A(net200),
    .B(clknet_1_1__leaf_net202),
    .C(net78),
    .X(net203));
 sky130_fd_sc_hd__and2_1 c226 (.A(net201),
    .B(net199),
    .X(net204));
 sky130_fd_sc_hd__and3_1 c227 (.A(net73),
    .B(net54),
    .C(net839),
    .X(net964));
 sky130_fd_sc_hd__and2_0 c228 (.A(net56),
    .B(net839),
    .X(net205));
 sky130_fd_sc_hd__and2_1 c229 (.A(net177),
    .B(net66),
    .X(net206));
 sky130_fd_sc_hd__a2111o_1 c230 (.A1(net154),
    .A2(net185),
    .B1(net50),
    .C1(net942),
    .D1(net989),
    .X(net207));
 sky130_fd_sc_hd__and3_1 c231 (.A(net205),
    .B(net206),
    .C(net839),
    .X(net208));
 sky130_fd_sc_hd__and2_1 c232 (.A(net157),
    .B(net1057),
    .X(net209));
 sky130_fd_sc_hd__and3_4 c233 (.A(net54),
    .B(net206),
    .C(net808),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_1 c234 (.A(net920),
    .X(net211));
 sky130_fd_sc_hd__a2111o_1 c235 (.A1(clknet_1_1__leaf_net197),
    .A2(net206),
    .B1(net154),
    .C1(net56),
    .D1(net210),
    .X(net212));
 sky130_fd_sc_hd__and2_0 c236 (.A(net210),
    .B(net808),
    .X(net213));
 sky130_fd_sc_hd__and3_1 c237 (.A(net206),
    .B(net209),
    .C(net210),
    .X(net214));
 sky130_fd_sc_hd__and3_1 c238 (.A(net43),
    .B(net191),
    .C(net213),
    .X(net215));
 sky130_fd_sc_hd__or4bb_2 c239 (.A(net211),
    .B(net213),
    .C_N(net989),
    .D_N(net71),
    .X(net216));
 sky130_fd_sc_hd__a2111o_1 c240 (.A1(net215),
    .A2(net205),
    .B1(net216),
    .C1(net43),
    .D1(clknet_1_0__leaf_net197),
    .X(net217));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(net209),
    .A1(net73),
    .A2(net215),
    .A3(net216),
    .S0(clknet_1_1__leaf_net217),
    .S1(net210),
    .X(net218));
 sky130_fd_sc_hd__and3_1 c242 (.A(net87),
    .B(clknet_1_0__leaf_net203),
    .C(net56),
    .X(net219));
 sky130_fd_sc_hd__and3_1 c243 (.A(net71),
    .B(net54),
    .C(net191),
    .X(net220));
 sky130_fd_sc_hd__or4bb_1 c244 (.A(net78),
    .B(net97),
    .C_N(net190),
    .D_N(net56),
    .X(net221));
 sky130_fd_sc_hd__or4bb_4 c245 (.A(net70),
    .B(net71),
    .C_N(net216),
    .D_N(net986),
    .X(net222));
 sky130_fd_sc_hd__buf_1 c246 (.A(net912),
    .X(net223));
 sky130_fd_sc_hd__mux4_1 c247 (.A0(net216),
    .A1(net89),
    .A2(net87),
    .A3(clknet_1_1__leaf_net977),
    .S0(net222),
    .S1(net1001),
    .X(net224));
 sky130_fd_sc_hd__and3_1 c248 (.A(net56),
    .B(net88),
    .C(net1001),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 c249 (.A(net912),
    .X(net226));
 sky130_fd_sc_hd__and2_1 c25 (.A(net944),
    .B(net948),
    .X(net0));
 sky130_fd_sc_hd__mux4_2 c250 (.A0(net66),
    .A1(net106),
    .A2(net210),
    .A3(net1001),
    .S0(net222),
    .S1(net101),
    .X(net976));
 sky130_fd_sc_hd__mux4_1 c251 (.A0(net67),
    .A1(net208),
    .A2(net216),
    .A3(net935),
    .S0(net191),
    .S1(net222),
    .X(net227));
 sky130_fd_sc_hd__and3_1 c252 (.A(net214),
    .B(net208),
    .C(net989),
    .X(net228));
 sky130_fd_sc_hd__mux4_1 c253 (.A0(net102),
    .A1(net222),
    .A2(net1001),
    .A3(clknet_1_1__leaf_net965),
    .S0(net990),
    .S1(net807),
    .X(net229));
 sky130_fd_sc_hd__buf_1 c254 (.A(net921),
    .X(net230));
 sky130_fd_sc_hd__and3_1 c255 (.A(clknet_1_1__leaf_net203),
    .B(net230),
    .C(net71),
    .X(net971));
 sky130_fd_sc_hd__mux4_1 c256 (.A0(net163),
    .A1(net230),
    .A2(clknet_1_1__leaf_net977),
    .A3(net222),
    .S0(net1001),
    .S1(clknet_1_1__leaf_net971),
    .X(net231));
 sky130_fd_sc_hd__and3_1 c257 (.A(net153),
    .B(net105),
    .C(net56),
    .X(net232));
 sky130_fd_sc_hd__mux4_1 c258 (.A0(net232),
    .A1(net228),
    .A2(clknet_1_1__leaf_net971),
    .A3(net222),
    .S0(net145),
    .S1(net1001),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_1 c259 (.A(net764),
    .X(net234));
 sky130_fd_sc_hd__and2_2 c26 (.A(net955),
    .B(net957),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c260 (.A0(net89),
    .A1(net106),
    .A2(net91),
    .A3(net70),
    .S0(net223),
    .S1(net785),
    .X(net235));
 sky130_fd_sc_hd__buf_2 c261 (.A(net929),
    .X(net236));
 sky130_fd_sc_hd__mux4_1 c262 (.A0(net106),
    .A1(net220),
    .A2(net230),
    .A3(net223),
    .S0(net236),
    .S1(net235),
    .X(net237));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net234),
    .A1(net235),
    .A2(net236),
    .A3(net785),
    .S0(net844),
    .S1(net848),
    .X(net238));
 sky130_fd_sc_hd__and2_1 c264 (.A(net941),
    .B(net119),
    .X(net239));
 sky130_fd_sc_hd__and2_0 c265 (.A(net956),
    .B(net997),
    .X(net240));
 sky130_fd_sc_hd__and2_1 c266 (.A(net240),
    .B(net997),
    .X(net241));
 sky130_fd_sc_hd__and2_2 c267 (.A(net240),
    .B(net116),
    .X(net242));
 sky130_fd_sc_hd__and3_2 c268 (.A(net111),
    .B(net935),
    .C(net240),
    .X(net243));
 sky130_fd_sc_hd__and3_4 c269 (.A(net943),
    .B(net242),
    .C(net123),
    .X(net244));
 sky130_fd_sc_hd__and3_1 c27 (.A(net947),
    .B(net951),
    .C(net950),
    .X(net2));
 sky130_fd_sc_hd__and3_4 c270 (.A(net121),
    .B(net239),
    .C(net243),
    .X(net245));
 sky130_fd_sc_hd__and2_1 c271 (.A(net979),
    .B(net243),
    .X(net246));
 sky130_fd_sc_hd__and3_1 c272 (.A(net123),
    .B(net127),
    .C(net116),
    .X(net247));
 sky130_fd_sc_hd__and3_1 c273 (.A(net112),
    .B(net242),
    .C(net243),
    .X(net248));
 sky130_fd_sc_hd__and2_0 c274 (.A(net239),
    .B(net954),
    .X(net249));
 sky130_fd_sc_hd__and2_1 c275 (.A(net246),
    .B(net126),
    .X(net250));
 sky130_fd_sc_hd__and2_1 c276 (.A(net249),
    .B(net125),
    .X(net251));
 sky130_fd_sc_hd__and3_1 c277 (.A(net249),
    .B(net248),
    .C(net251),
    .X(net252));
 sky130_fd_sc_hd__and2_0 c278 (.A(net241),
    .B(net243),
    .X(net253));
 sky130_fd_sc_hd__and2_1 c279 (.A(net248),
    .B(net956),
    .X(net254));
 sky130_fd_sc_hd__and2_4 c28 (.A(net1),
    .B(net2),
    .X(net3));
 sky130_fd_sc_hd__and2_1 c280 (.A(net251),
    .B(net254),
    .X(net255));
 sky130_fd_sc_hd__and3_2 c281 (.A(net248),
    .B(net245),
    .C(net243),
    .X(net256));
 sky130_fd_sc_hd__and3_1 c282 (.A(net247),
    .B(net126),
    .C(net256),
    .X(net257));
 sky130_fd_sc_hd__and3_1 c283 (.A(net252),
    .B(net256),
    .C(net257),
    .X(net258));
 sky130_fd_sc_hd__a2111o_2 c284 (.A1(net127),
    .A2(net248),
    .B1(net252),
    .C1(net255),
    .D1(net251),
    .X(net259));
 sky130_fd_sc_hd__or4bb_2 c285 (.A(net994),
    .B(net251),
    .C_N(net258),
    .D_N(net245),
    .X(net260));
 sky130_fd_sc_hd__and3_2 c286 (.A(net243),
    .B(net257),
    .C(net951),
    .X(net261));
 sky130_fd_sc_hd__and2_2 c287 (.A(net119),
    .B(net139),
    .X(net262));
 sky130_fd_sc_hd__buf_1 c288 (.A(clknet_1_0__leaf_net814),
    .X(net263));
 sky130_fd_sc_hd__and3_2 c289 (.A(net946),
    .B(net135),
    .C(net4),
    .X(net264));
 sky130_fd_sc_hd__mux4_2 c29 (.A0(net955),
    .A1(net3),
    .A2(net1),
    .A3(net944),
    .S0(net936),
    .S1(net950),
    .X(net4));
 sky130_fd_sc_hd__and2_1 c290 (.A(net257),
    .B(net993),
    .X(net265));
 sky130_fd_sc_hd__and3_1 c291 (.A(net265),
    .B(net993),
    .C(net832),
    .X(net266));
 sky130_fd_sc_hd__and2_1 c292 (.A(net136),
    .B(net266),
    .X(net267));
 sky130_fd_sc_hd__and3_1 c293 (.A(net7),
    .B(net261),
    .C(net832),
    .X(net268));
 sky130_fd_sc_hd__buf_1 c294 (.A(clknet_1_0__leaf_net814),
    .X(net269));
 sky130_fd_sc_hd__and2_2 c295 (.A(net260),
    .B(net833),
    .X(net270));
 sky130_fd_sc_hd__and3_2 c296 (.A(net266),
    .B(net270),
    .C(net18),
    .X(net271));
 sky130_fd_sc_hd__mux4_1 c297 (.A0(net0),
    .A1(net267),
    .A2(net270),
    .A3(net1059),
    .S0(net262),
    .S1(net993),
    .X(net272));
 sky130_fd_sc_hd__buf_1 c298 (.A(clknet_1_1__leaf_net924),
    .X(net273));
 sky130_fd_sc_hd__and3_1 c299 (.A(clknet_1_1__leaf_net273),
    .B(net241),
    .C(net270),
    .X(net274));
 sky130_fd_sc_hd__and2_1 c30 (.A(net4),
    .B(net3),
    .X(net5));
 sky130_fd_sc_hd__sdfrtp_1 c300 (.CLK(clknet_4_4_0_clk),
    .D(clknet_1_0__leaf_net274),
    .RESET_B(net271),
    .SCD(net950),
    .SCE(net851),
    .Q(net275));
 sky130_fd_sc_hd__or4bb_2 c301 (.A(net275),
    .B(net267),
    .C_N(net954),
    .D_N(net832),
    .X(net276));
 sky130_fd_sc_hd__and3_1 c302 (.A(net141),
    .B(net270),
    .C(net851),
    .X(net277));
 sky130_fd_sc_hd__buf_1 c303 (.A(net919),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_4 c304 (.A(net931),
    .X(net983));
 sky130_fd_sc_hd__mux4_1 c305 (.A0(net131),
    .A1(net275),
    .A2(net278),
    .A3(net256),
    .S0(net262),
    .S1(net243),
    .X(net279));
 sky130_fd_sc_hd__buf_1 c306 (.A(clknet_1_1__leaf_net922),
    .X(net280));
 sky130_fd_sc_hd__and3_1 c307 (.A(net278),
    .B(clknet_1_0__leaf_net273),
    .C(clknet_1_1__leaf_net814),
    .X(net281));
 sky130_fd_sc_hd__and2_0 c308 (.A(net139),
    .B(net245),
    .X(net282));
 sky130_fd_sc_hd__and3_1 c309 (.A(net260),
    .B(clknet_1_0__leaf_net172),
    .C(net21),
    .X(net283));
 sky130_fd_sc_hd__and2_1 c31 (.A(net2),
    .B(net943),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 c310 (.A(net737),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_2 c311 (.A(net737),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_1 c312 (.A(net794),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_1 c313 (.A(net794),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_1 c314 (.A(net931),
    .X(net288));
 sky130_fd_sc_hd__and2_1 c315 (.A(net29),
    .B(net165),
    .X(net968));
 sky130_fd_sc_hd__sdfbbn_1 c316 (.CLK_N(clknet_4_7_0_clk),
    .D(net284),
    .RESET_B(net995),
    .SCD(net285),
    .SCE(net955),
    .SET_B(net36),
    .Q(net290),
    .Q_N(net289));
 sky130_fd_sc_hd__and3_1 c317 (.A(net159),
    .B(clknet_1_0__leaf_net280),
    .C(net289),
    .X(net291));
 sky130_fd_sc_hd__buf_1 c318 (.A(clknet_1_0__leaf_net923),
    .X(net292));
 sky130_fd_sc_hd__and3_1 c319 (.A(net1058),
    .B(net268),
    .C(net992),
    .X(net293));
 sky130_fd_sc_hd__and3_2 c32 (.A(net3),
    .B(net958),
    .C(net5),
    .X(net7));
 sky130_fd_sc_hd__and3_1 c320 (.A(clknet_1_1__leaf_net172),
    .B(net285),
    .C(net287),
    .X(net294));
 sky130_fd_sc_hd__or4bb_1 c321 (.A(net292),
    .B(net290),
    .C_N(clknet_1_0__leaf_net294),
    .D_N(net992),
    .X(net295));
 sky130_fd_sc_hd__sdfbbn_2 c322 (.CLK_N(clknet_4_6_0_clk),
    .D(net286),
    .RESET_B(clknet_1_0__leaf_net294),
    .SCD(clknet_1_1__leaf_net295),
    .SCE(net992),
    .SET_B(net245),
    .Q(net960),
    .Q_N(net296));
 sky130_fd_sc_hd__buf_1 c323 (.A(net928),
    .X(net297));
 sky130_fd_sc_hd__a2111o_1 c324 (.A1(net139),
    .A2(net943),
    .B1(net992),
    .C1(net960),
    .D1(net156),
    .X(net298));
 sky130_fd_sc_hd__mux4_1 c325 (.A0(net166),
    .A1(net983),
    .A2(clknet_1_0__leaf_net295),
    .A3(net960),
    .S0(net285),
    .S1(net36),
    .X(net299));
 sky130_fd_sc_hd__mux4_1 c326 (.A0(net26),
    .A1(net261),
    .A2(clknet_1_0__leaf_net295),
    .A3(net992),
    .S0(net983),
    .S1(net852),
    .X(net300));
 sky130_fd_sc_hd__sdfbbp_1 c327 (.CLK(clknet_4_6_0_clk),
    .D(clknet_1_1__leaf_net295),
    .RESET_B(net286),
    .SCD(net170),
    .SCE(net852),
    .SET_B(net1013),
    .Q(net302),
    .Q_N(net301));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(net290),
    .A1(net979),
    .A2(net301),
    .A3(net794),
    .S0(net852),
    .S1(net853),
    .X(net303));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net303),
    .A1(net32),
    .A2(net302),
    .A3(net26),
    .S0(net296),
    .S1(net853),
    .X(net304));
 sky130_fd_sc_hd__and2_2 c33 (.A(net952),
    .B(net956),
    .X(net8));
 sky130_fd_sc_hd__buf_1 c330 (.X(net305));
 sky130_fd_sc_hd__buf_1 c331 (.A(net739),
    .X(net306));
 sky130_fd_sc_hd__buf_1 c332 (.A(clknet_1_1__leaf_net923),
    .X(net307));
 sky130_fd_sc_hd__and3_1 c333 (.A(net162),
    .B(net42),
    .C(net182),
    .X(net308));
 sky130_fd_sc_hd__mux4_1 c334 (.A0(net57),
    .A1(clknet_1_1__leaf_net965),
    .A2(net268),
    .A3(net306),
    .S0(net16),
    .S1(clknet_1_0__leaf_net842),
    .X(net309));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(net305),
    .A1(net32),
    .A2(net33),
    .A3(clknet_1_0__leaf_net842),
    .S0(clknet_1_0__leaf_net843),
    .S1(net854),
    .X(net310));
 sky130_fd_sc_hd__and2_0 c336 (.A(net794),
    .B(clknet_1_0__leaf_net841),
    .X(net311));
 sky130_fd_sc_hd__mux4_1 c337 (.A0(net36),
    .A1(net306),
    .A2(net960),
    .A3(clknet_1_0__leaf_net192),
    .S0(net305),
    .S1(clknet_1_1__leaf_net307),
    .X(net312));
 sky130_fd_sc_hd__and2_4 c338 (.A(net59),
    .B(net856),
    .X(net313));
 sky130_fd_sc_hd__a2111o_1 c339 (.A1(net313),
    .A2(net34),
    .B1(net42),
    .C1(clknet_1_1__leaf_net291),
    .D1(net854),
    .X(net314));
 sky130_fd_sc_hd__and3_1 c34 (.A(net5),
    .B(net949),
    .C(net2),
    .X(net9));
 sky130_fd_sc_hd__and2_0 c340 (.A(clknet_1_1__leaf_net294),
    .B(net855),
    .X(net315));
 sky130_fd_sc_hd__or4bb_1 c341 (.A(net311),
    .B(net57),
    .C_N(net992),
    .D_N(clknet_1_1__leaf_net307),
    .X(net316));
 sky130_fd_sc_hd__sdfsbp_1 c342 (.CLK(clknet_4_12_0_clk),
    .D(clknet_1_0__leaf_net291),
    .SCD(net1006),
    .SCE(net151),
    .SET_B(clknet_1_0__leaf_net310),
    .Q(net318),
    .Q_N(net317));
 sky130_fd_sc_hd__sdfbbn_1 c343 (.CLK_N(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net310),
    .RESET_B(net318),
    .SCD(net960),
    .SCE(clknet_1_1__leaf_net291),
    .SET_B(clknet_1_0__leaf_net192),
    .Q(net320),
    .Q_N(net319));
 sky130_fd_sc_hd__sdfbbn_1 c344 (.CLK_N(clknet_4_12_0_clk),
    .D(net16),
    .RESET_B(clknet_1_0__leaf_net316),
    .SCD(net317),
    .SCE(net3),
    .SET_B(clknet_1_1__leaf_net294),
    .Q(net322),
    .Q_N(net321));
 sky130_fd_sc_hd__and3_2 c345 (.A(net288),
    .B(net14),
    .C(net57),
    .X(net323));
 sky130_fd_sc_hd__mux4_1 c346 (.A0(clknet_1_1__leaf_net192),
    .A1(net306),
    .A2(net162),
    .A3(clknet_1_0__leaf_net280),
    .S0(net305),
    .S1(clknet_1_0__leaf_net841),
    .X(net324));
 sky130_fd_sc_hd__or4bb_1 c347 (.A(clknet_1_0__leaf_net315),
    .B(net33),
    .C_N(net185),
    .D_N(net986),
    .X(net325));
 sky130_fd_sc_hd__mux4_1 c348 (.A0(net308),
    .A1(net306),
    .A2(net323),
    .A3(clknet_1_1__leaf_net316),
    .S0(net42),
    .S1(clknet_1_0__leaf_net842),
    .X(net326));
 sky130_fd_sc_hd__buf_1 c349 (.A(clknet_1_0__leaf_net922),
    .X(net327));
 sky130_fd_sc_hd__and2_2 c35 (.A(net5),
    .B(net0),
    .X(net10));
 sky130_fd_sc_hd__and3_1 c350 (.A(clknet_1_1__leaf_net314),
    .B(net318),
    .C(net819),
    .X(net328));
 sky130_fd_sc_hd__sdfsbp_1 c351 (.CLK(clknet_4_12_0_clk),
    .D(net313),
    .SCD(net322),
    .SCE(clknet_1_1__leaf_net315),
    .SET_B(clknet_1_0__leaf_net327),
    .Q(net330),
    .Q_N(net329));
 sky130_fd_sc_hd__clkbuf_1 c352 (.A(net741),
    .X(net331));
 sky130_fd_sc_hd__and3_1 c353 (.A(net318),
    .B(net989),
    .C(net77),
    .X(net332));
 sky130_fd_sc_hd__buf_1 c354 (.A(net741),
    .X(net333));
 sky130_fd_sc_hd__sdfstp_1 c355 (.CLK(clknet_4_14_0_clk),
    .D(net32),
    .SCD(net84),
    .SCE(clknet_1_1__leaf_net218),
    .SET_B(net990),
    .Q(net334));
 sky130_fd_sc_hd__buf_1 c356 (.A(net748),
    .X(net335));
 sky130_fd_sc_hd__sdfbbp_1 c357 (.CLK(clknet_4_9_0_clk),
    .D(clknet_1_0__leaf_net316),
    .RESET_B(net335),
    .SCD(clknet_1_0__leaf_net328),
    .SCE(clknet_1_1__leaf_net842),
    .SET_B(net852),
    .Q(net337),
    .Q_N(net336));
 sky130_fd_sc_hd__clkbuf_2 c358 (.A(net747),
    .X(net338));
 sky130_fd_sc_hd__and2_0 c359 (.A(clknet_1_0__leaf_net202),
    .B(net321),
    .X(net339));
 sky130_fd_sc_hd__and3_1 c36 (.A(net948),
    .B(net5),
    .C(net10),
    .X(net11));
 sky130_fd_sc_hd__buf_1 c360 (.A(net759),
    .X(net340));
 sky130_fd_sc_hd__and2_0 c361 (.A(net335),
    .B(net338),
    .X(net341));
 sky130_fd_sc_hd__and3_1 c362 (.A(net73),
    .B(net990),
    .C(net857),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_1 c363 (.A(net759),
    .X(net343));
 sky130_fd_sc_hd__buf_1 c364 (.A(net765),
    .X(net344));
 sky130_fd_sc_hd__and3_1 c365 (.A(clknet_1_1__leaf_net212),
    .B(net329),
    .C(net333),
    .X(net345));
 sky130_fd_sc_hd__sdfstp_1 c366 (.CLK(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net274),
    .SCD(net338),
    .SCE(net990),
    .SET_B(net24),
    .Q(net346));
 sky130_fd_sc_hd__or4bb_1 c367 (.A(net343),
    .B(net276),
    .C_N(net346),
    .D_N(net994),
    .X(net347));
 sky130_fd_sc_hd__a2111o_1 c368 (.A1(net334),
    .A2(net343),
    .B1(net338),
    .C1(net936),
    .D1(clknet_1_1__leaf_net217),
    .X(net348));
 sky130_fd_sc_hd__a2111o_1 c369 (.A1(net330),
    .A2(clknet_1_0__leaf_net212),
    .B1(net344),
    .C1(net790),
    .D1(net852),
    .X(net962));
 sky130_fd_sc_hd__and2_1 c37 (.A(net11),
    .B(net1),
    .X(net12));
 sky130_fd_sc_hd__mux4_1 c370 (.A0(net331),
    .A1(clknet_1_1__leaf_net348),
    .A2(net318),
    .A3(net320),
    .S0(clknet_1_0__leaf_net962),
    .S1(net210),
    .X(net349));
 sky130_fd_sc_hd__sdfbbn_2 c371 (.CLK_N(clknet_4_14_0_clk),
    .D(net341),
    .RESET_B(net346),
    .SCD(clknet_1_0__leaf_net962),
    .SCE(net317),
    .SET_B(net994),
    .Q(net959),
    .Q_N(net350));
 sky130_fd_sc_hd__sdfbbn_1 c372 (.CLK_N(clknet_4_14_0_clk),
    .D(net342),
    .RESET_B(net1035),
    .SCD(net317),
    .SCE(clknet_1_0__leaf_net962),
    .SET_B(net858),
    .Q(net352),
    .Q_N(net351));
 sky130_fd_sc_hd__a2111o_1 c373 (.A1(net959),
    .A2(net351),
    .B1(clknet_1_1__leaf_net962),
    .C1(clknet_1_1__leaf_net842),
    .D1(net858),
    .X(net353));
 sky130_fd_sc_hd__mux4_1 c374 (.A0(net84),
    .A1(net236),
    .A2(net351),
    .A3(net987),
    .S0(net846),
    .S1(net1040),
    .X(net354));
 sky130_fd_sc_hd__a2111o_1 c375 (.A1(net941),
    .A2(net73),
    .B1(net338),
    .C1(net350),
    .D1(net807),
    .X(net355));
 sky130_fd_sc_hd__or4bb_1 c376 (.A(net97),
    .B(net1001),
    .C_N(net225),
    .D_N(net222),
    .X(net356));
 sky130_fd_sc_hd__a2111o_1 c377 (.A1(net210),
    .A2(clknet_1_0__leaf_net327),
    .B1(net338),
    .C1(net936),
    .D1(net845),
    .X(net357));
 sky130_fd_sc_hd__or4bb_4 c378 (.A(net939),
    .B(net84),
    .C_N(net146),
    .D_N(net352),
    .X(net358));
 sky130_fd_sc_hd__or4bb_4 c379 (.A(net88),
    .B(net63),
    .C_N(net358),
    .D_N(net807),
    .X(net967));
 sky130_fd_sc_hd__a2111o_1 c38 (.A1(net8),
    .A2(net944),
    .B1(net12),
    .C1(net936),
    .D1(net951),
    .X(net13));
 sky130_fd_sc_hd__mux4_1 c380 (.A0(net3),
    .A1(net994),
    .A2(net18),
    .A3(net358),
    .S0(clknet_1_0__leaf_net327),
    .S1(net852),
    .X(net359));
 sky130_fd_sc_hd__a2111o_1 c381 (.A1(net357),
    .A2(net225),
    .B1(net987),
    .C1(net358),
    .D1(net847),
    .X(net974));
 sky130_fd_sc_hd__or4bb_1 c382 (.A(net91),
    .B(net358),
    .C_N(clknet_1_1__leaf_net345),
    .D_N(net236),
    .X(net360));
 sky130_fd_sc_hd__a2111o_1 c383 (.A1(net222),
    .A2(net976),
    .B1(net1019),
    .C1(net967),
    .D1(net990),
    .X(net361));
 sky130_fd_sc_hd__or4bb_1 c384 (.A(net358),
    .B(net101),
    .C_N(net73),
    .D_N(net807),
    .X(net362));
 sky130_fd_sc_hd__mux4_1 c385 (.A0(net235),
    .A1(net987),
    .A2(net73),
    .A3(net358),
    .S0(net63),
    .S1(net1036),
    .X(net363));
 sky130_fd_sc_hd__sdfbbp_1 c386 (.CLK(clknet_4_14_0_clk),
    .D(clknet_1_0__leaf_net345),
    .RESET_B(net210),
    .SCD(net967),
    .SCE(net847),
    .SET_B(net852),
    .Q(net365),
    .Q_N(net364));
 sky130_fd_sc_hd__mux4_1 c387 (.A0(net359),
    .A1(net365),
    .A2(net362),
    .A3(net63),
    .S0(net338),
    .S1(net358),
    .X(net969));
 sky130_fd_sc_hd__or4bb_1 c388 (.A(net236),
    .B(net364),
    .C_N(net847),
    .D_N(net850),
    .X(net973));
 sky130_fd_sc_hd__mux4_1 c389 (.A0(net226),
    .A1(net362),
    .A2(net364),
    .A3(net786),
    .S0(net807),
    .S1(net859),
    .X(net366));
 sky130_fd_sc_hd__and2_4 c39 (.A(net12),
    .B(net13),
    .X(net14));
 sky130_fd_sc_hd__sdfbbn_1 c390 (.CLK_N(clknet_4_14_0_clk),
    .D(net354),
    .RESET_B(net356),
    .SCD(net365),
    .SCE(net1001),
    .SET_B(net236),
    .Q(net367));
 sky130_fd_sc_hd__mux4_2 c391 (.A0(net225),
    .A1(net1001),
    .A2(net210),
    .A3(net366),
    .S0(net967),
    .S1(net364),
    .X(net368));
 sky130_fd_sc_hd__mux4_1 c392 (.A0(net226),
    .A1(net338),
    .A2(net368),
    .A3(clknet_1_0__leaf_net969),
    .S0(clknet_1_0__leaf_net327),
    .S1(net101),
    .X(net369));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net366),
    .A1(net236),
    .A2(net368),
    .A3(net365),
    .S0(net1001),
    .S1(net296),
    .X(net370));
 sky130_fd_sc_hd__mux4_1 c394 (.A0(net101),
    .A1(net367),
    .A2(net358),
    .A3(net366),
    .S0(net222),
    .S1(net368),
    .X(net371));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net355),
    .A1(net358),
    .A2(clknet_1_1__leaf_net965),
    .A3(net368),
    .S0(net979),
    .S1(net859),
    .X(net372));
 sky130_fd_sc_hd__and2_0 c396 (.A(net129),
    .B(net258),
    .X(net373));
 sky130_fd_sc_hd__and2_2 c397 (.A(net260),
    .B(net112),
    .X(net374));
 sky130_fd_sc_hd__and2_1 c398 (.A(net126),
    .B(net254),
    .X(net375));
 sky130_fd_sc_hd__and2_2 c399 (.A(net957),
    .B(net242),
    .X(net376));
 sky130_fd_sc_hd__or4bb_2 c40 (.A(net11),
    .B(net937),
    .C_N(net9),
    .D_N(net14),
    .X(net15));
 sky130_fd_sc_hd__and2_1 c400 (.A(net375),
    .B(net120),
    .X(net377));
 sky130_fd_sc_hd__and2_0 c401 (.A(net247),
    .B(net375),
    .X(net378));
 sky130_fd_sc_hd__and2_2 c402 (.A(net373),
    .B(net256),
    .X(net379));
 sky130_fd_sc_hd__and2_1 c403 (.A(net122),
    .B(net253),
    .X(net380));
 sky130_fd_sc_hd__and2_2 c404 (.A(net938),
    .B(net379),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_1 c405 (.A(net723),
    .X(net382));
 sky130_fd_sc_hd__and2_4 c406 (.A(net254),
    .B(net375),
    .X(net383));
 sky130_fd_sc_hd__and2_0 c407 (.A(net255),
    .B(net379),
    .X(net384));
 sky130_fd_sc_hd__and2_1 c408 (.A(net379),
    .B(net382),
    .X(net385));
 sky130_fd_sc_hd__dlymetal6s2s_1 c409 (.A(net724),
    .X(net386));
 sky130_fd_sc_hd__a2111o_2 c41 (.A1(net15),
    .A2(net14),
    .B1(net955),
    .C1(net13),
    .D1(net11),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 c410 (.A(net933),
    .X(net387));
 sky130_fd_sc_hd__and3_1 c411 (.A(net382),
    .B(net255),
    .C(net379),
    .X(net388));
 sky130_fd_sc_hd__sdfbbn_1 c412 (.CLK_N(clknet_4_1_0_clk),
    .D(net388),
    .RESET_B(net1023),
    .SCD(net377),
    .SCE(net385),
    .SET_B(net383),
    .Q(net390),
    .Q_N(net389));
 sky130_fd_sc_hd__sdfstp_2 c413 (.CLK(clknet_4_1_0_clk),
    .D(net116),
    .SCD(net377),
    .SCE(net388),
    .SET_B(net383),
    .Q(net391));
 sky130_fd_sc_hd__or4bb_1 c414 (.A(net378),
    .B(net389),
    .C_N(net385),
    .D_N(net245),
    .X(net392));
 sky130_fd_sc_hd__sdfbbp_1 c415 (.CLK(clknet_4_1_0_clk),
    .D(net384),
    .RESET_B(net385),
    .SCD(net388),
    .SCE(net374),
    .SET_B(net1024),
    .Q(net394),
    .Q_N(net393));
 sky130_fd_sc_hd__a2111o_1 c416 (.A1(net393),
    .A2(net377),
    .B1(net389),
    .C1(net994),
    .D1(net795),
    .X(net395));
 sky130_fd_sc_hd__or4bb_1 c417 (.A(net394),
    .B(net390),
    .C_N(net384),
    .D_N(net386),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_1 c418 (.A(net736),
    .X(net397));
 sky130_fd_sc_hd__dlymetal6s2s_1 c419 (.A(net735),
    .X(net398));
 sky130_fd_sc_hd__or4bb_2 c42 (.A(net9),
    .B(net12),
    .C_N(net11),
    .D_N(net15),
    .X(net17));
 sky130_fd_sc_hd__and2_0 c420 (.A(net373),
    .B(net398),
    .X(net399));
 sky130_fd_sc_hd__and3_1 c421 (.A(net18),
    .B(clknet_1_0__leaf_net281),
    .C(net953),
    .X(net400));
 sky130_fd_sc_hd__and2_0 c422 (.A(net129),
    .B(net134),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_1 c423 (.A(net751),
    .X(net402));
 sky130_fd_sc_hd__and2_0 c424 (.A(net261),
    .B(net398),
    .X(net403));
 sky130_fd_sc_hd__and2_1 c425 (.A(net134),
    .B(net374),
    .X(net404));
 sky130_fd_sc_hd__and2_2 c426 (.A(net253),
    .B(net994),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_1 c427 (.A(net754),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_1 c428 (.A(net763),
    .X(net407));
 sky130_fd_sc_hd__and2_0 c429 (.A(net403),
    .B(net391),
    .X(net408));
 sky130_fd_sc_hd__mux4_2 c43 (.A0(net14),
    .A1(net13),
    .A2(net6),
    .A3(net9),
    .S0(net1),
    .S1(net10),
    .X(net18));
 sky130_fd_sc_hd__buf_1 c430 (.A(net761),
    .X(net409));
 sky130_fd_sc_hd__and2_2 c431 (.A(net399),
    .B(net991),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 c432 (.A0(net942),
    .A1(net991),
    .A2(net979),
    .A3(net398),
    .S0(clknet_1_0__leaf_net281),
    .S1(net993),
    .X(net411));
 sky130_fd_sc_hd__a2111o_1 c433 (.A1(clknet_1_0__leaf_net263),
    .A2(net380),
    .B1(net410),
    .C1(clknet_1_0__leaf_net411),
    .D1(net991),
    .X(net412));
 sky130_fd_sc_hd__or4bb_1 c434 (.A(net244),
    .B(net410),
    .C_N(net402),
    .X(net413));
 sky130_fd_sc_hd__mux4_1 c435 (.A0(net277),
    .A1(net253),
    .A2(net403),
    .A3(clknet_1_1__leaf_net263),
    .S0(net410),
    .S1(net979),
    .X(net414));
 sky130_fd_sc_hd__buf_1 c436 (.A(clknet_1_0__leaf_net924),
    .X(net415));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(clknet_1_0__leaf_net273),
    .A1(net270),
    .A2(clknet_1_0__leaf_net415),
    .A3(net410),
    .S0(net389),
    .S1(net381),
    .X(net416));
 sky130_fd_sc_hd__dlymetal6s2s_1 c438 (.A(net751),
    .X(net417));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net410),
    .A1(net398),
    .A2(net417),
    .A3(clknet_1_0__leaf_net415),
    .S0(net991),
    .S1(net865),
    .X(net418));
 sky130_fd_sc_hd__and2_0 c44 (.A(net950),
    .B(net952),
    .X(net19));
 sky130_fd_sc_hd__and2_0 c440 (.A(net133),
    .B(clknet_1_0__leaf_net415),
    .X(net419));
 sky130_fd_sc_hd__and2_0 c441 (.A(net390),
    .B(net14),
    .X(net420));
 sky130_fd_sc_hd__and2_0 c442 (.A(net420),
    .B(clknet_1_1__leaf_net411),
    .X(net421));
 sky130_fd_sc_hd__and2_0 c443 (.A(net995),
    .B(net865),
    .X(net422));
 sky130_fd_sc_hd__and2_0 c444 (.A(net376),
    .B(net992),
    .X(net423));
 sky130_fd_sc_hd__and2_0 c445 (.A(net124),
    .B(net285),
    .X(net424));
 sky130_fd_sc_hd__and3_2 c446 (.A(net406),
    .B(net960),
    .C(net995),
    .X(net425));
 sky130_fd_sc_hd__and3_1 c447 (.A(net421),
    .B(net245),
    .C(net995),
    .X(net426));
 sky130_fd_sc_hd__and3_1 c448 (.A(net285),
    .B(clknet_1_0__leaf_net294),
    .C(net293),
    .X(net427));
 sky130_fd_sc_hd__mux4_1 c449 (.A0(net282),
    .A1(net951),
    .A2(net301),
    .A3(net285),
    .S0(net383),
    .S1(net823),
    .X(net428));
 sky130_fd_sc_hd__and2_1 c45 (.A(net40),
    .B(net8),
    .X(net20));
 sky130_fd_sc_hd__and2_1 c450 (.A(net424),
    .B(net397),
    .X(net429));
 sky130_fd_sc_hd__mux4_1 c451 (.A0(clknet_1_1__leaf_net281),
    .A1(net995),
    .A2(net936),
    .A3(net297),
    .S0(net285),
    .S1(net997),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_1 c452 (.A(net932),
    .X(net431));
 sky130_fd_sc_hd__and3_2 c453 (.A(net951),
    .B(net150),
    .C(net820),
    .X(net432));
 sky130_fd_sc_hd__mux4_1 c454 (.A0(net419),
    .A1(net431),
    .A2(net432),
    .A3(net425),
    .S0(clknet_1_0__leaf_net427),
    .S1(net261),
    .X(net433));
 sky130_fd_sc_hd__mux4_1 c455 (.A0(net398),
    .A1(net133),
    .A2(net21),
    .A3(net432),
    .S0(clknet_1_0__leaf_net427),
    .S1(net1003),
    .X(net434));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(net431),
    .A1(net409),
    .A2(net1006),
    .A3(net398),
    .S0(net864),
    .S1(net1004),
    .X(net435));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(clknet_1_0__leaf_net411),
    .A1(net435),
    .A2(net993),
    .A3(clknet_1_1__leaf_net427),
    .S0(net432),
    .S1(net1003),
    .X(net436));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(net397),
    .A1(net432),
    .A2(net995),
    .A3(clknet_1_1__leaf_net427),
    .S0(net1004),
    .S1(net870),
    .X(net437));
 sky130_fd_sc_hd__a2111o_1 c459 (.A1(net432),
    .A2(net425),
    .B1(net823),
    .C1(net1003),
    .D1(net870),
    .X(net438));
 sky130_fd_sc_hd__and2_4 c46 (.A(net949),
    .B(net8),
    .X(net21));
 sky130_fd_sc_hd__mux4_2 c460 (.A0(net435),
    .A1(net438),
    .A2(net425),
    .A3(net432),
    .S0(net1004),
    .S1(net870),
    .X(net439));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net438),
    .A1(net250),
    .A2(net439),
    .A3(net151),
    .S0(net1004),
    .S1(net870),
    .X(net440));
 sky130_fd_sc_hd__a2111o_1 c462 (.A1(net187),
    .A2(net439),
    .B1(clknet_1_0__leaf_net307),
    .C1(net979),
    .D1(net991),
    .X(net441));
 sky130_fd_sc_hd__and3_1 c463 (.A(net270),
    .B(net187),
    .C(net183),
    .X(net442));
 sky130_fd_sc_hd__and3_1 c464 (.A(net409),
    .B(clknet_1_1__leaf_net327),
    .C(net986),
    .X(net443));
 sky130_fd_sc_hd__mux4_1 c465 (.A0(net442),
    .A1(clknet_1_1__leaf_net427),
    .A2(net183),
    .A3(net439),
    .S0(net245),
    .S1(net986),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_2 c466 (.A(net916),
    .X(net978));
 sky130_fd_sc_hd__sedfxbp_1 c467 (.CLK(clknet_4_9_0_clk),
    .D(net271),
    .DE(net186),
    .SCD(net936),
    .SCE(net870),
    .Q(net446),
    .Q_N(net445));
 sky130_fd_sc_hd__clkbuf_1 c468 (.A(net915),
    .X(net447));
 sky130_fd_sc_hd__and3_1 c469 (.A(net429),
    .B(net322),
    .C(net991),
    .X(net448));
 sky130_fd_sc_hd__and2_1 c47 (.A(net2),
    .B(net16),
    .X(net22));
 sky130_fd_sc_hd__a2111o_1 c470 (.A1(net1007),
    .A2(net978),
    .B1(clknet_1_0__leaf_net307),
    .C1(net818),
    .D1(net870),
    .X(net449));
 sky130_fd_sc_hd__and3_1 c471 (.A(net449),
    .B(net445),
    .C(net1003),
    .X(net450));
 sky130_fd_sc_hd__or4bb_1 c472 (.A(net151),
    .B(clknet_1_1__leaf_net307),
    .C_N(net994),
    .D_N(net1003),
    .X(net451));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(net268),
    .A1(clknet_1_1__leaf_net427),
    .A2(net439),
    .A3(net1006),
    .S0(clknet_1_1__leaf_net450),
    .S1(net1003),
    .X(net452));
 sky130_fd_sc_hd__and3_1 c474 (.A(net443),
    .B(net391),
    .C(net379),
    .X(net453));
 sky130_fd_sc_hd__mux4_1 c475 (.A0(net270),
    .A1(net439),
    .A2(clknet_1_1__leaf_net450),
    .A3(clknet_1_0__leaf_net453),
    .S0(net991),
    .S1(net820),
    .X(net454));
 sky130_fd_sc_hd__sedfxbp_1 c476 (.CLK(clknet_4_6_0_clk),
    .D(clknet_1_0__leaf_net307),
    .DE(clknet_1_0__leaf_net453),
    .SCD(net296),
    .SCE(net783),
    .Q(net455));
 sky130_fd_sc_hd__mux4_1 c477 (.A0(clknet_1_0__leaf_net307),
    .A1(clknet_1_1__leaf_net294),
    .A2(clknet_1_0__leaf_net451),
    .A3(clknet_1_0__leaf_net328),
    .S0(clknet_1_1__leaf_net450),
    .S1(net111),
    .X(net456));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(net430),
    .A1(net1009),
    .A2(clknet_1_1__leaf_net314),
    .A3(clknet_1_0__leaf_net453),
    .S0(net296),
    .S1(net955),
    .X(net457));
 sky130_fd_sc_hd__sedfxtp_4 c479 (.CLK(clknet_4_6_0_clk),
    .D(net245),
    .DE(clknet_1_0__leaf_net451),
    .SCD(clknet_1_0__leaf_net453),
    .SCE(net1008),
    .Q(net458));
 sky130_fd_sc_hd__and2_0 c48 (.A(net20),
    .B(net19),
    .X(net23));
 sky130_fd_sc_hd__or4bb_1 c480 (.A(net1021),
    .B(net42),
    .C_N(net439),
    .D_N(net1003),
    .X(net459));
 sky130_fd_sc_hd__and3_1 c481 (.A(net379),
    .B(clknet_1_1__leaf_net294),
    .C(clknet_1_1__leaf_net450),
    .X(net460));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(net447),
    .A1(clknet_1_0__leaf_net460),
    .A2(clknet_1_1__leaf_net450),
    .A3(net458),
    .S0(net1008),
    .S1(clknet_1_1__leaf_net453),
    .X(net461));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net1008),
    .A1(clknet_1_0__leaf_net460),
    .A2(net321),
    .A3(clknet_1_1__leaf_net450),
    .S0(net871),
    .S1(net872),
    .X(net462));
 sky130_fd_sc_hd__and3_1 c484 (.A(clknet_1_1__leaf_net328),
    .B(clknet_1_0__leaf_net217),
    .C(net1002),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_1 c485 (.A(net911),
    .X(net464));
 sky130_fd_sc_hd__a2111o_1 c486 (.A1(clknet_1_0__leaf_net316),
    .A2(clknet_1_0__leaf_net328),
    .B1(net986),
    .C1(clknet_1_0__leaf_net962),
    .D1(net63),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_1 c487 (.A(net911),
    .X(net466));
 sky130_fd_sc_hd__and3_1 c488 (.A(net380),
    .B(net466),
    .C(net63),
    .X(net467));
 sky130_fd_sc_hd__and3_1 c489 (.A(net466),
    .B(net987),
    .C(net993),
    .X(net970));
 sky130_fd_sc_hd__and2_4 c49 (.A(net938),
    .B(net21),
    .X(net24));
 sky130_fd_sc_hd__and3_2 c490 (.A(net337),
    .B(net446),
    .C(net868),
    .X(net980));
 sky130_fd_sc_hd__and3_2 c491 (.A(net996),
    .B(net793),
    .C(net868),
    .X(net468));
 sky130_fd_sc_hd__and3_1 c492 (.A(net322),
    .B(net84),
    .C(net980),
    .X(net469));
 sky130_fd_sc_hd__and3_1 c493 (.A(net344),
    .B(net970),
    .C(net350),
    .X(net470));
 sky130_fd_sc_hd__and3_1 c494 (.A(net111),
    .B(net24),
    .C(net336),
    .X(net471));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(net470),
    .A1(net469),
    .A2(clknet_1_1__leaf_net453),
    .A3(net1006),
    .S0(net335),
    .S1(net868),
    .X(net472));
 sky130_fd_sc_hd__mux4_2 c496 (.A0(net446),
    .A1(net970),
    .A2(clknet_1_1__leaf_net328),
    .A3(net978),
    .S0(net980),
    .S1(net1004),
    .X(net473));
 sky130_fd_sc_hd__and3_1 c497 (.A(clknet_1_1__leaf_net451),
    .B(net471),
    .C(net829),
    .X(net474));
 sky130_fd_sc_hd__and3_1 c498 (.A(net448),
    .B(net471),
    .C(net871),
    .X(net475));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(net959),
    .A1(clknet_1_1__leaf_net962),
    .A2(net984),
    .A3(clknet_1_1__leaf_net453),
    .S0(net789),
    .S1(net874),
    .X(net476));
 sky130_fd_sc_hd__and2_1 c50 (.A(net12),
    .B(net21),
    .X(net25));
 sky130_fd_sc_hd__a2111o_1 c500 (.A1(clknet_1_0__leaf_net217),
    .A2(net344),
    .B1(net18),
    .C1(net445),
    .D1(net876),
    .X(net477));
 sky130_fd_sc_hd__and3_1 c501 (.A(net993),
    .B(net980),
    .C(net875),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(clknet_1_1__leaf_net453),
    .A1(net467),
    .A2(net939),
    .A3(net478),
    .S0(net968),
    .S1(net996),
    .X(net479));
 sky130_fd_sc_hd__sdfbbn_1 c503 (.CLK_N(clknet_4_11_0_clk),
    .D(net463),
    .RESET_B(net478),
    .SCD(net471),
    .SCE(net84),
    .SET_B(net876),
    .Q(net481),
    .Q_N(net480));
 sky130_fd_sc_hd__and3_1 c504 (.A(net475),
    .B(net471),
    .C(net481),
    .X(net482));
 sky130_fd_sc_hd__and3_1 c505 (.A(net464),
    .B(net474),
    .C(net875),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c509 (.A0(net937),
    .A1(clknet_1_0__leaf_net473),
    .A2(net480),
    .A3(clknet_1_0__leaf_net971),
    .S0(clknet_1_0__leaf_net327),
    .S1(clknet_1_0__leaf_net863),
    .X(net484));
 sky130_fd_sc_hd__and2_2 c51 (.A(net22),
    .B(net25),
    .X(net26));
 sky130_fd_sc_hd__a2111o_1 c510 (.A1(clknet_1_1__leaf_net327),
    .A2(net480),
    .B1(net146),
    .C1(clknet_1_0__leaf_net863),
    .D1(net874),
    .X(net485));
 sky130_fd_sc_hd__a2111o_1 c511 (.A1(net146),
    .A2(clknet_1_1__leaf_net327),
    .B1(net860),
    .C1(net861),
    .D1(net877),
    .X(net486));
 sky130_fd_sc_hd__sdfbbn_1 c512 (.CLK_N(clknet_4_11_0_clk),
    .D(net950),
    .RESET_B(clknet_1_1__leaf_net473),
    .SCD(net1038),
    .SCE(net983),
    .SET_B(clknet_1_0__leaf_net862),
    .Q(net488),
    .Q_N(net487));
 sky130_fd_sc_hd__a2111o_1 c513 (.A1(net63),
    .A2(net125),
    .B1(net996),
    .C1(net115),
    .D1(net487),
    .X(net489));
 sky130_fd_sc_hd__or4bb_1 c514 (.A(net489),
    .B(net488),
    .C_N(net980),
    .D_N(net845),
    .X(net490));
 sky130_fd_sc_hd__a2111o_1 c515 (.A1(net352),
    .A2(net488),
    .B1(net983),
    .C1(net989),
    .D1(clknet_1_1__leaf_net327),
    .X(net491));
 sky130_fd_sc_hd__a2111o_1 c516 (.A1(net486),
    .A2(clknet_1_1__leaf_net451),
    .B1(net488),
    .C1(net1006),
    .D1(net989),
    .X(net492));
 sky130_fd_sc_hd__a2111o_1 c517 (.A1(net492),
    .A2(net481),
    .B1(net487),
    .C1(net860),
    .D1(clknet_1_1__leaf_net862),
    .X(net493));
 sky130_fd_sc_hd__a2111o_1 c518 (.A1(net362),
    .A2(clknet_1_1__leaf_net491),
    .B1(clknet_1_1__leaf_net327),
    .C1(net487),
    .D1(net860),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c519 (.A0(net221),
    .A1(net989),
    .A2(net950),
    .A3(net987),
    .S0(clknet_1_1__leaf_net863),
    .S1(net878),
    .X(net495));
 sky130_fd_sc_hd__and2_2 c52 (.A(net19),
    .B(net25),
    .X(net27));
 sky130_fd_sc_hd__mux4_1 c520 (.A0(net244),
    .A1(net368),
    .A2(net488),
    .A3(clknet_1_1__leaf_net451),
    .S0(net350),
    .S1(net849),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c521 (.A0(clknet_1_0__leaf_net485),
    .A1(clknet_1_0__leaf_net491),
    .A2(net967),
    .A3(net488),
    .S0(net871),
    .S1(net879),
    .X(net497));
 sky130_fd_sc_hd__a2111o_1 c522 (.A1(net481),
    .A2(net495),
    .B1(clknet_1_1__leaf_net485),
    .C1(clknet_1_1__leaf_net327),
    .D1(net1012),
    .X(net498));
 sky130_fd_sc_hd__a2111o_1 c523 (.A1(net115),
    .A2(net488),
    .B1(clknet_1_0__leaf_net497),
    .C1(net980),
    .D1(net1012),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c524 (.A0(net490),
    .A1(clknet_1_1__leaf_net497),
    .A2(net487),
    .A3(net978),
    .S0(net805),
    .S1(net1012),
    .X(net500));
 sky130_fd_sc_hd__sdfbbp_1 c525 (.CLK(clknet_4_11_0_clk),
    .D(net368),
    .RESET_B(clknet_1_0__leaf_net971),
    .SCD(net976),
    .SCE(net1039),
    .SET_B(net1012),
    .Q(net502),
    .Q_N(net501));
 sky130_fd_sc_hd__mux4_1 c526 (.A0(clknet_1_1__leaf_net327),
    .A1(net493),
    .A2(net502),
    .A3(net989),
    .S0(net487),
    .S1(net879),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c527 (.A0(net123),
    .A1(net494),
    .A2(net503),
    .A3(net501),
    .S0(net828),
    .S1(net879),
    .X(net504));
 sky130_fd_sc_hd__and2_0 c528 (.A(net246),
    .B(net250),
    .X(net505));
 sky130_fd_sc_hd__and2_1 c529 (.A(net390),
    .B(net374),
    .X(net506));
 sky130_fd_sc_hd__and2_0 c53 (.A(net23),
    .B(net40),
    .X(net28));
 sky130_fd_sc_hd__and2_0 c530 (.A(net505),
    .B(net374),
    .X(net507));
 sky130_fd_sc_hd__buf_1 c531 (.A(net831),
    .X(net508));
 sky130_fd_sc_hd__and3_1 c532 (.A(net375),
    .B(net942),
    .C(net795),
    .X(net509));
 sky130_fd_sc_hd__and2_0 c533 (.A(net387),
    .B(net383),
    .X(net510));
 sky130_fd_sc_hd__dlymetal6s2s_1 c534 (.A(net831),
    .X(net511));
 sky130_fd_sc_hd__and2_2 c535 (.A(net510),
    .B(net256),
    .X(net512));
 sky130_fd_sc_hd__clkbuf_1 c536 (.A(net750),
    .X(net513));
 sky130_fd_sc_hd__and2_2 c537 (.A(net509),
    .B(net117),
    .X(net514));
 sky130_fd_sc_hd__and2_0 c538 (.A(net395),
    .B(net511),
    .X(net515));
 sky130_fd_sc_hd__and2_1 c539 (.A(net511),
    .B(net386),
    .X(net516));
 sky130_fd_sc_hd__and2_1 c54 (.A(net25),
    .B(net0),
    .X(net29));
 sky130_fd_sc_hd__or4bb_2 c540 (.A(net515),
    .B(net510),
    .C_N(net514),
    .D_N(net997),
    .X(net517));
 sky130_fd_sc_hd__or4bb_1 c541 (.A(net512),
    .B(net244),
    .C_N(net509),
    .D_N(net513),
    .X(net518));
 sky130_fd_sc_hd__and2_1 c542 (.A(net508),
    .B(net518),
    .X(net519));
 sky130_fd_sc_hd__and2_0 c543 (.A(net518),
    .B(net508),
    .X(net520));
 sky130_fd_sc_hd__and2_0 c544 (.A(net519),
    .B(net515),
    .X(net521));
 sky130_fd_sc_hd__or4bb_2 c545 (.A(net258),
    .B(net519),
    .C_N(net514),
    .D_N(net511),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 c546 (.A0(net516),
    .A1(net519),
    .A2(net521),
    .A3(net511),
    .S0(net508),
    .S1(net514),
    .X(net523));
 sky130_fd_sc_hd__and2_1 c547 (.A(net511),
    .B(net812),
    .X(net524));
 sky130_fd_sc_hd__mux4_1 c548 (.A0(net521),
    .A1(net519),
    .A2(net395),
    .A3(net524),
    .S0(net514),
    .S1(net516),
    .X(net525));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(net516),
    .A1(net520),
    .A2(net508),
    .A3(net511),
    .S0(net519),
    .S1(net812),
    .X(net526));
 sky130_fd_sc_hd__and2_0 c55 (.A(net23),
    .B(net22),
    .X(net30));
 sky130_fd_sc_hd__and2_0 c550 (.A(net265),
    .B(net517),
    .X(net527));
 sky130_fd_sc_hd__and2_1 c551 (.A(net401),
    .B(net376),
    .X(net528));
 sky130_fd_sc_hd__and2_0 c552 (.A(net250),
    .B(net994),
    .X(net529));
 sky130_fd_sc_hd__clkbuf_1 c553 (.A(net816),
    .X(net530));
 sky130_fd_sc_hd__and2_0 c554 (.A(net524),
    .B(net528),
    .X(net531));
 sky130_fd_sc_hd__sedfxtp_4 c555 (.CLK(clknet_4_1_0_clk),
    .D(net531),
    .DE(net949),
    .SCD(net528),
    .SCE(net991),
    .Q(net532));
 sky130_fd_sc_hd__and2_4 c556 (.A(net528),
    .B(net866),
    .X(net533));
 sky130_fd_sc_hd__clkbuf_1 c557 (.A(net926),
    .X(net534));
 sky130_fd_sc_hd__and2_0 c558 (.A(net534),
    .B(net524),
    .X(net535));
 sky130_fd_sc_hd__and2_0 c559 (.A(clknet_1_0__leaf_net269),
    .B(net417),
    .X(net536));
 sky130_fd_sc_hd__and2_1 c56 (.A(net28),
    .B(net23),
    .X(net31));
 sky130_fd_sc_hd__and2_0 c560 (.A(net536),
    .B(net528),
    .X(net537));
 sky130_fd_sc_hd__buf_1 c561 (.A(net816),
    .X(net538));
 sky130_fd_sc_hd__and2_0 c562 (.A(net528),
    .B(net867),
    .X(net539));
 sky130_fd_sc_hd__buf_1 c563 (.A(net750),
    .X(net540));
 sky130_fd_sc_hd__and2_0 c564 (.A(net513),
    .B(net417),
    .X(net541));
 sky130_fd_sc_hd__clkbuf_1 c565 (.A(net761),
    .X(net542));
 sky130_fd_sc_hd__buf_2 c566 (.A(net762),
    .X(net543));
 sky130_fd_sc_hd__buf_1 c567 (.A(net925),
    .X(net544));
 sky130_fd_sc_hd__mux4_1 c568 (.A0(net417),
    .A1(net544),
    .A2(net534),
    .A3(net541),
    .S0(clknet_1_1__leaf_net537),
    .S1(net533),
    .X(net545));
 sky130_fd_sc_hd__and3_4 c569 (.A(net542),
    .B(net544),
    .C(net529),
    .X(net546));
 sky130_fd_sc_hd__and3_2 c57 (.A(net30),
    .B(net20),
    .C(net31),
    .X(net32));
 sky130_fd_sc_hd__and2_1 c570 (.A(net514),
    .B(net546),
    .X(net547));
 sky130_fd_sc_hd__clkbuf_4 c571 (.A(net754),
    .X(net548));
 sky130_fd_sc_hd__and3_2 c572 (.A(net517),
    .B(net949),
    .C(net1004),
    .X(net549));
 sky130_fd_sc_hd__clkbuf_2 c573 (.A(net732),
    .X(net550));
 sky130_fd_sc_hd__mux4_1 c574 (.A0(net440),
    .A1(net423),
    .A2(net1),
    .A3(net993),
    .S0(net550),
    .S1(net992),
    .X(net551));
 sky130_fd_sc_hd__buf_1 c575 (.A(net732),
    .X(net552));
 sky130_fd_sc_hd__and3_1 c576 (.A(net426),
    .B(net547),
    .C(net134),
    .X(net553));
 sky130_fd_sc_hd__and3_1 c577 (.A(net544),
    .B(net823),
    .C(net1004),
    .X(net554));
 sky130_fd_sc_hd__and3_1 c578 (.A(net538),
    .B(net549),
    .C(clknet_1_1__leaf_net415),
    .X(net555));
 sky130_fd_sc_hd__and3_2 c579 (.A(net293),
    .B(net997),
    .C(net817),
    .X(net556));
 sky130_fd_sc_hd__and2_2 c58 (.A(net27),
    .B(net28),
    .X(net33));
 sky130_fd_sc_hd__and2_0 c580 (.A(net425),
    .B(net817),
    .X(net557));
 sky130_fd_sc_hd__and2_0 c581 (.A(net557),
    .B(net514),
    .X(net558));
 sky130_fd_sc_hd__and2_2 c582 (.A(net554),
    .B(net1004),
    .X(net559));
 sky130_fd_sc_hd__and3_1 c583 (.A(net374),
    .B(net261),
    .C(net558),
    .X(net560));
 sky130_fd_sc_hd__and3_1 c584 (.A(net297),
    .B(net517),
    .C(net559),
    .X(net561));
 sky130_fd_sc_hd__mux4_1 c585 (.A0(net111),
    .A1(net561),
    .A2(net1000),
    .A3(net548),
    .S0(net995),
    .S1(net1018),
    .X(net562));
 sky130_fd_sc_hd__sedfxtp_2 c586 (.CLK(clknet_4_3_0_clk),
    .D(net547),
    .DE(net517),
    .SCD(clknet_1_0__leaf_net977),
    .SCE(net556),
    .Q(net563));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(net995),
    .A1(net562),
    .A2(net563),
    .A3(clknet_1_1__leaf_net553),
    .S0(net543),
    .S1(net870),
    .X(net564));
 sky130_fd_sc_hd__sdfrbp_1 c588 (.CLK(clknet_4_3_0_clk),
    .D(net561),
    .RESET_B(net562),
    .SCD(net563),
    .SCE(net559),
    .Q(net566),
    .Q_N(net565));
 sky130_fd_sc_hd__a2111o_1 c589 (.A1(net561),
    .A2(net565),
    .B1(net514),
    .C1(net820),
    .D1(net880),
    .X(net567));
 sky130_fd_sc_hd__and3_2 c59 (.A(net31),
    .B(net15),
    .C(net33),
    .X(net34));
 sky130_fd_sc_hd__a2111o_1 c590 (.A1(net1),
    .A2(net556),
    .B1(net550),
    .C1(net566),
    .D1(net560),
    .X(net568));
 sky130_fd_sc_hd__clkbuf_1 c591 (.A(net1028),
    .X(net569));
 sky130_fd_sc_hd__a2111o_1 c592 (.A1(net558),
    .A2(net1052),
    .B1(net425),
    .C1(net569),
    .D1(net556),
    .X(net570));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(net560),
    .A1(net569),
    .A2(net563),
    .A3(net546),
    .S0(net1),
    .S1(net880),
    .X(net571));
 sky130_fd_sc_hd__mux4_1 c594 (.A0(clknet_1_0__leaf_net314),
    .A1(net183),
    .A2(net242),
    .A3(clknet_1_0__leaf_net965),
    .S0(net548),
    .S1(net556),
    .X(net572));
 sky130_fd_sc_hd__sdfbbn_1 c595 (.CLK_N(clknet_4_3_0_clk),
    .D(net540),
    .RESET_B(net323),
    .SCD(clknet_1_1__leaf_net555),
    .SCE(net301),
    .SET_B(net556),
    .Q(net574),
    .Q_N(net573));
 sky130_fd_sc_hd__mux4_2 c596 (.A0(net543),
    .A1(net566),
    .A2(net14),
    .A3(net991),
    .S0(net559),
    .S1(net784),
    .X(net575));
 sky130_fd_sc_hd__or4bb_1 c597 (.A(net991),
    .B(net39),
    .C_N(net559),
    .D_N(net543),
    .X(net576));
 sky130_fd_sc_hd__sdfbbn_1 c598 (.CLK_N(clknet_4_3_0_clk),
    .D(net323),
    .RESET_B(net950),
    .SCD(net458),
    .SCE(net988),
    .SET_B(net1000),
    .Q(net578),
    .Q_N(net577));
 sky130_fd_sc_hd__mux4_1 c599 (.A0(net559),
    .A1(net42),
    .A2(clknet_1_0__leaf_net450),
    .A3(net988),
    .S0(net870),
    .S1(net1002),
    .X(net579));
 sky130_fd_sc_hd__and3_1 c60 (.A(net40),
    .B(net949),
    .C(net30),
    .X(net35));
 sky130_fd_sc_hd__a2111o_1 c600 (.A1(net242),
    .A2(clknet_1_0__leaf_net314),
    .B1(net42),
    .C1(net984),
    .D1(net872),
    .X(net580));
 sky130_fd_sc_hd__mux4_1 c601 (.A0(net579),
    .A1(net566),
    .A2(net242),
    .A3(net533),
    .S0(net182),
    .S1(net546),
    .X(net581));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(clknet_1_0__leaf_net555),
    .A1(net994),
    .A2(net988),
    .A3(clknet_1_0__leaf_net450),
    .S0(net459),
    .S1(clknet_1_0__leaf_net963),
    .X(net582));
 sky130_fd_sc_hd__or4bb_1 c603 (.A(net183),
    .B(net578),
    .C_N(net988),
    .D_N(clknet_1_0__leaf_net883),
    .X(net583));
 sky130_fd_sc_hd__a2111o_1 c604 (.A1(clknet_1_0__leaf_net450),
    .A2(clknet_1_0__leaf_net583),
    .B1(net405),
    .C1(net988),
    .D1(clknet_1_0__leaf_net883),
    .X(net961));
 sky130_fd_sc_hd__a2111o_1 c605 (.A1(clknet_1_0__leaf_net583),
    .A2(net988),
    .B1(net546),
    .C1(net577),
    .D1(clknet_1_0__leaf_net883),
    .X(net584));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net422),
    .A1(net993),
    .A2(net1006),
    .A3(clknet_1_0__leaf_net961),
    .S0(net135),
    .S1(net1000),
    .X(net585));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(net323),
    .A1(clknet_1_0__leaf_net584),
    .A2(net42),
    .A3(net391),
    .S0(clknet_1_0__leaf_net961),
    .S1(clknet_1_0__leaf_net882),
    .X(net586));
 sky130_fd_sc_hd__or4bb_1 c608 (.A(clknet_1_1__leaf_net584),
    .B(clknet_1_0__leaf_net450),
    .C_N(clknet_1_1__leaf_net883),
    .D_N(net885),
    .X(net587));
 sky130_fd_sc_hd__mux4_1 c609 (.A0(clknet_1_0__leaf_net584),
    .A1(net988),
    .A2(clknet_1_0__leaf_net587),
    .A3(net810),
    .S0(clknet_1_1__leaf_net882),
    .S1(net885),
    .X(net588));
 sky130_fd_sc_hd__and3_2 c61 (.A(net35),
    .B(net34),
    .C(net33),
    .X(net36));
 sky130_fd_sc_hd__a2111o_1 c610 (.A1(net540),
    .A2(clknet_1_1__leaf_net583),
    .B1(net182),
    .C1(net811),
    .D1(net887),
    .X(net982));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(clknet_1_1__leaf_net982),
    .A1(net988),
    .A2(clknet_1_0__leaf_net961),
    .A3(clknet_1_1__leaf_net584),
    .S0(net872),
    .S1(clknet_1_1__leaf_net883),
    .X(net589));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(net42),
    .A1(clknet_1_1__leaf_net587),
    .A2(clknet_1_1__leaf_net982),
    .A3(clknet_1_1__leaf_net961),
    .S0(net872),
    .S1(net886),
    .X(net590));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(net556),
    .A1(clknet_1_0__leaf_net982),
    .A2(clknet_1_0__leaf_net587),
    .A3(clknet_1_0__leaf_net965),
    .S0(net884),
    .S1(net889),
    .X(net591));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(net546),
    .A1(net585),
    .A2(clknet_1_1__leaf_net982),
    .A3(clknet_1_0__leaf_net589),
    .S0(net884),
    .S1(net888),
    .X(net592));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(clknet_1_1__leaf_net587),
    .A1(net405),
    .A2(net549),
    .A3(net821),
    .S0(net888),
    .S1(net890),
    .X(net593));
 sky130_fd_sc_hd__a2111o_1 c616 (.A1(net340),
    .A2(net468),
    .B1(net993),
    .C1(net1000),
    .D1(net1006),
    .X(net594));
 sky130_fd_sc_hd__a2111o_1 c617 (.A1(net477),
    .A2(net978),
    .B1(net996),
    .C1(net264),
    .D1(net881),
    .X(net595));
 sky130_fd_sc_hd__or4bb_1 c618 (.A(net559),
    .B(net575),
    .C_N(net543),
    .D_N(net873),
    .X(net596));
 sky130_fd_sc_hd__or4bb_1 c619 (.A(net549),
    .B(net596),
    .C_N(clknet_1_0__leaf_net962),
    .D_N(net1002),
    .X(net597));
 sky130_fd_sc_hd__mux4_1 c62 (.A0(net22),
    .A1(net28),
    .A2(net25),
    .A3(net34),
    .S0(net27),
    .S1(net14),
    .X(net37));
 sky130_fd_sc_hd__or4bb_2 c620 (.A(net543),
    .B(net1000),
    .C_N(net468),
    .D_N(net559),
    .X(net966));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(net996),
    .A1(clknet_1_0__leaf_net962),
    .A2(net988),
    .A3(net800),
    .S0(net1004),
    .S1(net891),
    .X(net598));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(clknet_1_1__leaf_net460),
    .A1(net468),
    .A2(net1006),
    .A3(net350),
    .S0(net543),
    .S1(net892),
    .X(net599));
 sky130_fd_sc_hd__a2111o_1 c623 (.A1(clknet_1_0__leaf_net589),
    .A2(net134),
    .B1(net549),
    .C1(net1004),
    .D1(clknet_1_1__leaf_net963),
    .X(net600));
 sky130_fd_sc_hd__sdfbbp_1 c624 (.CLK(clknet_4_11_0_clk),
    .D(net936),
    .RESET_B(net204),
    .SCD(net983),
    .SCE(net972),
    .SET_B(net892),
    .Q(net601));
 sky130_fd_sc_hd__sdfrbp_2 c625 (.CLK(clknet_4_10_0_clk),
    .D(net533),
    .RESET_B(net1029),
    .SCD(net1033),
    .SCE(clknet_1_1__leaf_net963),
    .Q(net603),
    .Q_N(net602));
 sky130_fd_sc_hd__a2111o_1 c626 (.A1(net302),
    .A2(clknet_1_1__leaf_net441),
    .B1(net24),
    .C1(net983),
    .D1(net891),
    .X(net604));
 sky130_fd_sc_hd__sdfbbn_1 c627 (.CLK_N(clknet_4_10_0_clk),
    .D(net204),
    .RESET_B(net601),
    .SCD(net966),
    .SCE(net603),
    .SET_B(net549),
    .Q(net606),
    .Q_N(net605));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net332),
    .A1(net574),
    .A2(net606),
    .A3(net602),
    .S0(net264),
    .S1(net1005),
    .X(net607));
 sky130_fd_sc_hd__a2111o_1 c629 (.A1(net988),
    .A2(net594),
    .B1(net302),
    .C1(net966),
    .D1(net602),
    .X(net608));
 sky130_fd_sc_hd__mux4_1 c63 (.A0(net19),
    .A1(net946),
    .A2(net35),
    .A3(net36),
    .S0(net31),
    .S1(net21),
    .X(net38));
 sky130_fd_sc_hd__sdfbbn_1 c630 (.CLK_N(clknet_4_9_0_clk),
    .D(net14),
    .RESET_B(clknet_1_1__leaf_net589),
    .SCD(net1000),
    .SCE(net543),
    .SET_B(net1002),
    .Q(net609));
 sky130_fd_sc_hd__mux4_2 c631 (.A0(net383),
    .A1(net970),
    .A2(net512),
    .A3(net602),
    .S0(net296),
    .S1(net605),
    .X(net610));
 sky130_fd_sc_hd__a2111o_1 c632 (.A1(net608),
    .A2(clknet_1_1__leaf_net589),
    .B1(net610),
    .C1(net891),
    .D1(net892),
    .X(net611));
 sky130_fd_sc_hd__sdfbbp_1 c633 (.CLK(clknet_4_11_0_clk),
    .D(net984),
    .RESET_B(clknet_1_0__leaf_net217),
    .SCD(net610),
    .SCE(clknet_1_1__leaf_net961),
    .SET_B(net989),
    .Q(net612));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net607),
    .A1(net980),
    .A2(net610),
    .A3(net966),
    .S0(net605),
    .S1(net829),
    .X(net613));
 sky130_fd_sc_hd__sdfbbn_1 c635 (.CLK_N(clknet_4_8_0_clk),
    .D(net1022),
    .RESET_B(net604),
    .SCD(net512),
    .SCE(net992),
    .SET_B(net605),
    .Q(net615),
    .Q_N(net614));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net612),
    .A1(net614),
    .A2(net966),
    .A3(net602),
    .S0(net1046),
    .S1(net893),
    .X(net616));
 sky130_fd_sc_hd__sdfbbn_1 c637 (.CLK_N(clknet_4_10_0_clk),
    .D(net610),
    .RESET_B(net616),
    .SCD(net1045),
    .SCE(net980),
    .SET_B(net1032),
    .Q(net618),
    .Q_N(net617));
 sky130_fd_sc_hd__and3_4 c64 (.A(net30),
    .B(net35),
    .C(net1051),
    .X(net39));
 sky130_fd_sc_hd__and2_1 c65 (.A(net954),
    .B(net1),
    .X(net40));
 sky130_fd_sc_hd__buf_1 c66 (.A(net804),
    .X(net41));
 sky130_fd_sc_hd__buf_1 c660 (.A(net803),
    .X(net619));
 sky130_fd_sc_hd__buf_1 c661 (.A(net803),
    .X(net620));
 sky130_fd_sc_hd__and2_0 c662 (.A(net239),
    .B(net110),
    .X(net621));
 sky130_fd_sc_hd__buf_1 c663 (.A(net802),
    .X(net622));
 sky130_fd_sc_hd__and2_1 c664 (.A(net620),
    .B(net120),
    .X(net623));
 sky130_fd_sc_hd__and2_1 c665 (.A(net120),
    .B(net622),
    .X(net624));
 sky130_fd_sc_hd__buf_1 c666 (.A(net802),
    .X(net625));
 sky130_fd_sc_hd__and2_2 c667 (.A(net621),
    .B(net375),
    .X(net626));
 sky130_fd_sc_hd__and2_0 c668 (.A(net520),
    .B(net626),
    .X(net627));
 sky130_fd_sc_hd__and2_0 c669 (.A(net376),
    .B(net624),
    .X(net628));
 sky130_fd_sc_hd__and2_2 c67 (.A(net948),
    .B(net27),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 c670 (.A(net830),
    .X(net629));
 sky130_fd_sc_hd__and2_1 c671 (.A(net391),
    .B(net386),
    .X(net630));
 sky130_fd_sc_hd__clkbuf_1 c672 (.A(net932),
    .X(net631));
 sky130_fd_sc_hd__and2_2 c673 (.A(net935),
    .B(net621),
    .X(net632));
 sky130_fd_sc_hd__and3_1 c674 (.A(net630),
    .B(net631),
    .C(net998),
    .X(net633));
 sky130_fd_sc_hd__and2_1 c675 (.A(net631),
    .B(net624),
    .X(net634));
 sky130_fd_sc_hd__clkbuf_1 c676 (.A(net830),
    .X(net635));
 sky130_fd_sc_hd__and3_1 c677 (.A(net632),
    .B(net998),
    .C(net633),
    .X(net636));
 sky130_fd_sc_hd__and3_1 c678 (.A(net628),
    .B(net620),
    .C(net633),
    .X(net637));
 sky130_fd_sc_hd__a2111o_1 c679 (.A1(net637),
    .A2(net632),
    .B1(net633),
    .C1(net628),
    .D1(net998),
    .X(net638));
 sky130_fd_sc_hd__and2_1 c68 (.A(net946),
    .B(net41),
    .X(net43));
 sky130_fd_sc_hd__a2111o_1 c680 (.A1(net633),
    .A2(net630),
    .B1(net638),
    .C1(net637),
    .D1(net998),
    .X(net639));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(net638),
    .A1(net636),
    .A2(net635),
    .A3(net619),
    .S0(net633),
    .S1(net998),
    .X(net640));
 sky130_fd_sc_hd__sdfrtn_1 c682 (.CLK_N(clknet_4_0_0_clk),
    .D(net1031),
    .RESET_B(net639),
    .SCD(net548),
    .SCE(clknet_1_0__leaf_net537),
    .Q(net641));
 sky130_fd_sc_hd__clkbuf_1 c683 (.A(net913),
    .X(net642));
 sky130_fd_sc_hd__dlymetal6s2s_1 c684 (.A(net913),
    .X(net643));
 sky130_fd_sc_hd__sdfrtp_4 c685 (.CLK(clknet_4_0_0_clk),
    .D(net386),
    .RESET_B(net522),
    .SCD(net532),
    .SCE(net643),
    .Q(net644));
 sky130_fd_sc_hd__clkbuf_1 c686 (.A(net934),
    .X(net645));
 sky130_fd_sc_hd__buf_1 c687 (.A(net822),
    .X(net646));
 sky130_fd_sc_hd__and3_1 c688 (.A(net645),
    .B(net640),
    .C(net950),
    .X(net647));
 sky130_fd_sc_hd__and3_1 c689 (.A(net642),
    .B(clknet_1_0__leaf_net537),
    .C(net641),
    .X(net648));
 sky130_fd_sc_hd__and2_1 c69 (.A(net9),
    .B(net31),
    .X(net44));
 sky130_fd_sc_hd__and3_1 c690 (.A(net639),
    .B(net135),
    .C(net386),
    .X(net649));
 sky130_fd_sc_hd__clkbuf_1 c691 (.A(net822),
    .X(net650));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(net506),
    .A1(net244),
    .A2(net622),
    .A3(net636),
    .S0(net532),
    .S1(net546),
    .X(net651));
 sky130_fd_sc_hd__a2111o_1 c693 (.A1(net256),
    .A2(net533),
    .B1(net1026),
    .C1(net1056),
    .D1(net1014),
    .X(net652));
 sky130_fd_sc_hd__and3_1 c694 (.A(net650),
    .B(net623),
    .C(net383),
    .X(net653));
 sky130_fd_sc_hd__clkbuf_1 c695 (.A(net934),
    .X(net654));
 sky130_fd_sc_hd__and3_1 c696 (.A(net654),
    .B(net125),
    .C(net1047),
    .X(net655));
 sky130_fd_sc_hd__a2111o_1 c697 (.A1(net548),
    .A2(net625),
    .B1(net641),
    .C1(net532),
    .D1(net796),
    .X(net656));
 sky130_fd_sc_hd__and3_2 c698 (.A(net643),
    .B(net653),
    .C(net894),
    .X(net657));
 sky130_fd_sc_hd__and3_1 c699 (.A(net119),
    .B(net635),
    .C(net894),
    .X(net658));
 sky130_fd_sc_hd__and2_1 c70 (.A(net950),
    .B(net4),
    .X(net45));
 sky130_fd_sc_hd__and3_1 c700 (.A(net653),
    .B(net658),
    .C(net256),
    .X(net659));
 sky130_fd_sc_hd__buf_1 c701 (.A(net933),
    .X(net660));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net659),
    .A1(net548),
    .A2(net643),
    .A3(net998),
    .S0(net645),
    .S1(net634),
    .X(net661));
 sky130_fd_sc_hd__and3_1 c703 (.A(net660),
    .B(net661),
    .C(net659),
    .X(net662));
 sky130_fd_sc_hd__sdfbbp_1 c704 (.CLK(clknet_4_2_0_clk),
    .D(clknet_1_0__leaf_net553),
    .RESET_B(net999),
    .SCD(net244),
    .SCE(net662),
    .SET_B(net1020),
    .Q(net664),
    .Q_N(net663));
 sky130_fd_sc_hd__a2111o_1 c705 (.A1(net640),
    .A2(net551),
    .B1(net797),
    .C1(net1054),
    .D1(net1047),
    .X(net665));
 sky130_fd_sc_hd__a2111o_1 c706 (.A1(net655),
    .A2(net432),
    .B1(net550),
    .C1(clknet_1_0__leaf_net977),
    .D1(net1047),
    .X(net666));
 sky130_fd_sc_hd__buf_1 c707 (.A(net917),
    .X(net667));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(net425),
    .A1(net641),
    .A2(net546),
    .A3(net550),
    .S0(net999),
    .S1(net799),
    .X(net668));
 sky130_fd_sc_hd__and3_1 c709 (.A(net623),
    .B(net640),
    .C(net668),
    .X(net669));
 sky130_fd_sc_hd__and2_0 c71 (.A(net24),
    .B(net8),
    .X(net46));
 sky130_fd_sc_hd__and3_1 c710 (.A(net668),
    .B(net432),
    .C(net798),
    .X(net670));
 sky130_fd_sc_hd__and3_1 c711 (.A(net667),
    .B(net548),
    .C(net641),
    .X(net671));
 sky130_fd_sc_hd__a2111o_1 c712 (.A1(net649),
    .A2(net383),
    .B1(net376),
    .C1(net644),
    .D1(net998),
    .X(net672));
 sky130_fd_sc_hd__and3_1 c713 (.A(net636),
    .B(net662),
    .C(net644),
    .X(net673));
 sky130_fd_sc_hd__and3_1 c714 (.A(net641),
    .B(net626),
    .C(net425),
    .X(net674));
 sky130_fd_sc_hd__sdfbbn_1 c715 (.CLK_N(clknet_4_2_0_clk),
    .D(net673),
    .RESET_B(net667),
    .SCD(net670),
    .SCE(net432),
    .SET_B(net792),
    .Q(net676),
    .Q_N(net675));
 sky130_fd_sc_hd__and3_2 c716 (.A(net432),
    .B(net674),
    .C(net425),
    .X(net677));
 sky130_fd_sc_hd__a2111o_1 c717 (.A1(net953),
    .A2(net677),
    .B1(net998),
    .C1(net798),
    .D1(net1003),
    .X(net678));
 sky130_fd_sc_hd__a2111o_1 c718 (.A1(net550),
    .A2(net634),
    .B1(net667),
    .C1(net677),
    .D1(net880),
    .X(net679));
 sky130_fd_sc_hd__mux4_2 c719 (.A0(net656),
    .A1(net939),
    .A2(net676),
    .A3(net383),
    .S0(net677),
    .S1(net999),
    .X(net680));
 sky130_fd_sc_hd__and2_0 c72 (.A(net43),
    .B(net31),
    .X(net47));
 sky130_fd_sc_hd__a2111o_1 c720 (.A1(net939),
    .A2(net677),
    .B1(net985),
    .C1(net799),
    .D1(net880),
    .X(net681));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net679),
    .A1(net677),
    .A2(net681),
    .A3(net641),
    .S0(net985),
    .S1(net1048),
    .X(net682));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net622),
    .A1(net678),
    .A2(net669),
    .A3(net677),
    .S0(net985),
    .S1(net681),
    .X(net683));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net677),
    .A1(net681),
    .A2(net985),
    .A3(net548),
    .S0(net675),
    .S1(net1034),
    .X(net684));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net985),
    .A1(net677),
    .A2(net827),
    .A3(net894),
    .S0(net896),
    .S1(net897),
    .X(net685));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net671),
    .A1(net685),
    .A2(net677),
    .A3(net985),
    .S0(net797),
    .S1(net880),
    .X(net686));
 sky130_fd_sc_hd__or4bb_1 c726 (.A(net999),
    .B(net549),
    .C_N(net669),
    .D_N(net575),
    .X(net687));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net459),
    .A1(net1020),
    .A2(net135),
    .A3(net115),
    .S0(net1002),
    .S1(net890),
    .X(net688));
 sky130_fd_sc_hd__or4bb_1 c728 (.A(net664),
    .B(net670),
    .C_N(net657),
    .D_N(net881),
    .X(net689));
 sky130_fd_sc_hd__a2111o_1 c729 (.A1(net24),
    .A2(net1000),
    .B1(net18),
    .C1(net663),
    .D1(net244),
    .X(net690));
 sky130_fd_sc_hd__and2_0 c73 (.A(net6),
    .B(net37),
    .X(net48));
 sky130_fd_sc_hd__a2111o_1 c730 (.A1(net634),
    .A2(net672),
    .B1(net552),
    .C1(net458),
    .D1(net1005),
    .X(net691));
 sky130_fd_sc_hd__sdfrtp_1 c731 (.CLK(clknet_4_2_0_clk),
    .D(net646),
    .RESET_B(net688),
    .SCD(net657),
    .SCE(net985),
    .Q(net692));
 sky130_fd_sc_hd__or4bb_4 c732 (.A(net458),
    .B(net692),
    .C_N(net664),
    .D_N(net672),
    .X(net693));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(clknet_1_1__leaf_net456),
    .A1(net693),
    .A2(net672),
    .A3(net657),
    .S0(net1000),
    .S1(net868),
    .X(net694));
 sky130_fd_sc_hd__or4bb_1 c734 (.A(net1000),
    .B(net692),
    .C_N(clknet_1_0__leaf_net965),
    .D_N(net693),
    .X(net695));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net690),
    .A1(net692),
    .A2(net985),
    .A3(net657),
    .S0(net675),
    .S1(net632),
    .X(net696));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(net687),
    .A1(net670),
    .A2(net18),
    .A3(net24),
    .S0(net890),
    .S1(net1015),
    .X(net697));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net135),
    .A1(net548),
    .A2(net626),
    .A3(clknet_1_0__leaf_net441),
    .S0(net1000),
    .S1(net900),
    .X(net698));
 sky130_fd_sc_hd__mux4_2 c738 (.A0(net632),
    .A1(net646),
    .A2(net957),
    .A3(net693),
    .S0(net787),
    .S1(net881),
    .X(net699));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(net696),
    .A1(net634),
    .A2(clknet_1_0__leaf_net698),
    .A3(net699),
    .S0(net244),
    .S1(clknet_1_0__leaf_net456),
    .X(net700));
 sky130_fd_sc_hd__and2_1 c74 (.A(net37),
    .B(net44),
    .X(net49));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(net644),
    .A1(net681),
    .A2(net699),
    .A3(net985),
    .S0(net546),
    .S1(net899),
    .X(net701));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(clknet_1_0__leaf_net441),
    .A1(net699),
    .A2(net39),
    .A3(net881),
    .S0(net890),
    .S1(net901),
    .X(net702));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(net691),
    .A1(net644),
    .A2(net999),
    .A3(clknet_1_0__leaf_net965),
    .S0(net828),
    .S1(net901),
    .X(net703));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(net669),
    .A1(net942),
    .A2(net646),
    .A3(net699),
    .S0(net825),
    .S1(net901),
    .X(net704));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(net693),
    .A1(net699),
    .A2(net632),
    .A3(net1005),
    .S0(net901),
    .S1(net903),
    .X(net705));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(clknet_1_1__leaf_net698),
    .A1(net699),
    .A2(net383),
    .A3(net548),
    .S0(net787),
    .S1(net890),
    .X(net706));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net689),
    .A1(net699),
    .A2(net1005),
    .A3(net900),
    .S0(net901),
    .S1(clknet_1_0__leaf_net904),
    .X(net707));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(net676),
    .A1(net548),
    .A2(net826),
    .A3(net902),
    .S0(clknet_1_0__leaf_net904),
    .S1(net906),
    .X(net708));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net333),
    .A1(net618),
    .A2(net950),
    .A3(net793),
    .S0(net1002),
    .S1(net899),
    .X(net709));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net657),
    .A1(net709),
    .A2(net693),
    .A3(net533),
    .S0(net468),
    .S1(net899),
    .X(net710));
 sky130_fd_sc_hd__and2_2 c75 (.A(net48),
    .B(net41),
    .X(net50));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(net482),
    .A1(net575),
    .A2(net606),
    .A3(net603),
    .S0(net1005),
    .S1(net889),
    .X(net711));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net468),
    .A1(net693),
    .A2(net615),
    .A3(net617),
    .S0(net603),
    .S1(net994),
    .X(net712));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net603),
    .A1(net259),
    .A2(clknet_1_1__leaf_net977),
    .A3(clknet_1_0__leaf_net708),
    .S0(net1002),
    .S1(net901),
    .X(net713));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net676),
    .A1(net957),
    .A2(clknet_1_1__leaf_net441),
    .A3(net573),
    .S0(net806),
    .S1(net1002),
    .X(net714));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net339),
    .A1(net996),
    .A2(net985),
    .A3(net573),
    .S0(net657),
    .S1(net889),
    .X(net715));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net626),
    .A1(net483),
    .A2(net575),
    .A3(net996),
    .S0(net1002),
    .S1(net901),
    .X(net716));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net574),
    .A1(net711),
    .A2(clknet_1_1__leaf_net708),
    .A3(net615),
    .S0(net24),
    .S1(net603),
    .X(net717));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net533),
    .A1(net715),
    .A2(net614),
    .A3(clknet_1_0__leaf_net965),
    .S0(net895),
    .S1(clknet_1_1__leaf_net904),
    .X(net718));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net123),
    .A1(net881),
    .A2(net901),
    .A3(net906),
    .S0(net907),
    .S1(net908),
    .X(net719));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net712),
    .A1(net714),
    .A2(net716),
    .A3(clknet_1_0__leaf_net708),
    .S0(net693),
    .S1(net908),
    .X(net720));
 sky130_fd_sc_hd__and2_1 c76 (.A(net41),
    .B(net49),
    .X(net51));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net680),
    .A1(net806),
    .A2(net896),
    .A3(net905),
    .S0(net909),
    .S1(net910),
    .X(net721));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net719),
    .A1(net721),
    .A2(net996),
    .A3(net533),
    .S0(net1030),
    .S1(net910),
    .X(net722));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net606),
    .A1(net18),
    .A2(net680),
    .A3(net824),
    .S0(net909),
    .S1(net910));
 sky130_fd_sc_hd__clkbuf_1 c77 (.A(net804),
    .X(net52));
 sky130_fd_sc_hd__and2_1 c78 (.A(net45),
    .B(net49),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 c79 (.A(net804),
    .X(net54));
 sky130_fd_sc_hd__buf_1 c80 (.A(net749),
    .X(net55));
 sky130_fd_sc_hd__buf_2 c81 (.A(net749),
    .X(net56));
 sky130_fd_sc_hd__and2_2 c82 (.A(net37),
    .B(net55),
    .X(net57));
 sky130_fd_sc_hd__buf_1 c83 (.A(net930),
    .X(net58));
 sky130_fd_sc_hd__and2_4 c84 (.A(net52),
    .B(net834),
    .X(net59));
 sky130_fd_sc_hd__mux4_1 c85 (.A0(net10),
    .A1(net48),
    .A2(net44),
    .A3(net53),
    .S0(net41),
    .S1(net59),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 c86 (.A(net775),
    .X(net61));
 sky130_fd_sc_hd__mux4_1 c87 (.A0(net61),
    .A1(net34),
    .A2(net56),
    .A3(net53),
    .S0(net57),
    .S1(net1044),
    .X(net62));
 sky130_fd_sc_hd__and2_4 c88 (.A(net953),
    .B(net20),
    .X(net63));
 sky130_fd_sc_hd__and2_1 c89 (.A(net47),
    .B(net54),
    .X(net64));
 sky130_fd_sc_hd__sdfbbn_1 c90 (.CLK_N(clknet_4_13_0_clk),
    .D(net20),
    .RESET_B(net64),
    .SCD(net50),
    .SCE(net63),
    .SET_B(net838),
    .Q(net66),
    .Q_N(net65));
 sky130_fd_sc_hd__and2_1 c91 (.A(net1049),
    .B(net54),
    .X(net67));
 sky130_fd_sc_hd__and2_0 c92 (.A(net33),
    .B(net54),
    .X(net68));
 sky130_fd_sc_hd__and2_0 c93 (.A(net937),
    .B(net67),
    .X(net69));
 sky130_fd_sc_hd__and2_1 c94 (.A(net936),
    .B(net67),
    .X(net70));
 sky130_fd_sc_hd__and2_2 c95 (.A(net46),
    .B(net56),
    .X(net71));
 sky130_fd_sc_hd__and2_0 c96 (.A(net68),
    .B(net836),
    .X(net72));
 sky130_fd_sc_hd__and2_2 c97 (.A(net18),
    .B(net67),
    .X(net73));
 sky130_fd_sc_hd__and2_1 c98 (.A(net32),
    .B(net8),
    .X(net74));
 sky130_fd_sc_hd__and3_2 c99 (.A(net69),
    .B(net63),
    .C(net70),
    .X(net75));
 sky130_fd_sc_hd__sdfbbn_1 merge763 (.CLK_N(clknet_4_1_0_clk),
    .D(net385),
    .RESET_B(net383),
    .SCD(net377),
    .SCE(net381),
    .SET_B(net376),
    .Q(net724),
    .Q_N(net723));
 sky130_fd_sc_hd__mux4_1 merge764 (.A0(clknet_1_0__leaf_net348),
    .A1(net340),
    .A2(clknet_1_1__leaf_net280),
    .A3(clknet_1_1__leaf_net460),
    .S0(net1003),
    .S1(net1002),
    .X(net725));
 sky130_fd_sc_hd__mux4_1 merge765 (.A0(net190),
    .A1(net214),
    .A2(clknet_1_1__leaf_net977),
    .A3(net93),
    .S0(net63),
    .S1(net67),
    .X(net726));
 sky130_fd_sc_hd__or4bb_1 merge766 (.A(net47),
    .B(net51),
    .C_N(net52),
    .D_N(net53),
    .X(net727));
 sky130_fd_sc_hd__mux4_1 merge767 (.A0(net532),
    .A1(net623),
    .A2(net522),
    .A3(net935),
    .S0(net642),
    .S1(clknet_1_0__leaf_net537),
    .X(net728));
 sky130_fd_sc_hd__or4bb_1 merge768 (.A(net110),
    .B(net522),
    .C_N(net375),
    .D_N(net526),
    .X(net729));
 sky130_fd_sc_hd__sdfbbp_1 merge769 (.CLK(clknet_4_5_0_clk),
    .D(net143),
    .RESET_B(net150),
    .SCD(net156),
    .SCE(net112),
    .SET_B(net32),
    .Q(net731),
    .Q_N(net730));
 sky130_fd_sc_hd__sdfrtp_1 merge770 (.CLK(clknet_4_3_0_clk),
    .D(net304),
    .RESET_B(clknet_1_1__leaf_net415),
    .SCD(net547),
    .SCE(net1003),
    .Q(net732));
 sky130_fd_sc_hd__mux4_1 merge771 (.A0(net34),
    .A1(net54),
    .A2(net156),
    .A3(net51),
    .S0(net986),
    .S1(net840),
    .X(net733));
 sky130_fd_sc_hd__a2111o_1 merge772 (.A1(net50),
    .A2(net99),
    .B1(net3),
    .C1(net97),
    .D1(net74),
    .X(net734));
 sky130_fd_sc_hd__sdfsbp_1 merge773 (.CLK(clknet_4_4_0_clk),
    .D(net262),
    .SCD(net265),
    .SCE(net943),
    .SET_B(net271),
    .Q(net736),
    .Q_N(net735));
 sky130_fd_sc_hd__clkbuf_1 merge774 (.A(net919),
    .X(net737));
 sky130_fd_sc_hd__sdfbbn_1 merge775 (.CLK_N(clknet_4_7_0_clk),
    .RESET_B(net184),
    .SCD(net156),
    .SCE(net111),
    .SET_B(clknet_1_0__leaf_net841),
    .Q(net739),
    .Q_N(net305));
 sky130_fd_sc_hd__mux4_1 merge776 (.A0(net439),
    .A1(net39),
    .A2(net1008),
    .A3(net112),
    .S0(net391),
    .S1(net323),
    .X(net740));
 sky130_fd_sc_hd__buf_1 merge777 (.A(net822),
    .X(net741));
 sky130_fd_sc_hd__or4bb_1 merge778 (.A(net388),
    .B(net246),
    .C_N(net117),
    .D_N(net381),
    .X(net742));
 sky130_fd_sc_hd__or4bb_1 merge779 (.A(net21),
    .B(net74),
    .C_N(net82),
    .D_N(net81),
    .X(net743));
 sky130_fd_sc_hd__or4bb_1 merge780 (.A(net381),
    .B(net514),
    .C_N(net529),
    .D_N(clknet_1_1__leaf_net537),
    .X(net744));
 sky130_fd_sc_hd__or4bb_1 merge781 (.A(net81),
    .B(net67),
    .C_N(net199),
    .D_N(net154),
    .X(net745));
 sky130_fd_sc_hd__or4bb_1 merge782 (.A(net262),
    .B(net241),
    .C_N(net267),
    .D_N(net938),
    .X(net746));
 sky130_fd_sc_hd__sdfsbp_1 merge783 (.CLK(clknet_4_12_0_clk),
    .D(net198),
    .SCD(clknet_1_0__leaf_net218),
    .SCE(net33),
    .SET_B(clknet_1_1__leaf_net316),
    .Q(net748),
    .Q_N(net747));
 sky130_fd_sc_hd__clkbuf_1 merge784 (.A(net776),
    .X(net749));
 sky130_fd_sc_hd__sdfstp_1 merge785 (.CLK(clknet_4_1_0_clk),
    .D(net535),
    .SCD(net404),
    .SCE(net507),
    .SET_B(net511),
    .Q(net750));
 sky130_fd_sc_hd__sdfstp_1 merge786 (.CLK(clknet_4_1_0_clk),
    .D(net400),
    .SCD(net262),
    .SCE(net410),
    .SET_B(net809),
    .Q(net751));
 sky130_fd_sc_hd__or4bb_1 merge787 (.A(net278),
    .B(net156),
    .C_N(net283),
    .D_N(net271),
    .X(net752));
 sky130_fd_sc_hd__mux4_1 merge788 (.A0(net567),
    .A1(net563),
    .A2(net565),
    .A3(net551),
    .S0(net546),
    .S1(net533),
    .X(net753));
 sky130_fd_sc_hd__sdfstp_1 merge789 (.CLK(clknet_4_1_0_clk),
    .D(net241),
    .SCD(net262),
    .SCE(net404),
    .SET_B(net546),
    .Q(net754));
 sky130_fd_sc_hd__mux4_1 merge790 (.A0(net136),
    .A1(net262),
    .A2(clknet_1_0__leaf_net274),
    .A3(net36),
    .S0(net242),
    .S1(net170),
    .X(net755));
 sky130_fd_sc_hd__mux4_1 merge791 (.A0(net31),
    .A1(net33),
    .A2(net39),
    .A3(net169),
    .S0(net156),
    .S1(clknet_1_1__leaf_net813),
    .X(net756));
 sky130_fd_sc_hd__mux4_1 merge792 (.A0(net175),
    .A1(net50),
    .A2(net169),
    .A3(net73),
    .S0(net210),
    .S1(net1042),
    .X(net757));
 sky130_fd_sc_hd__mux4_1 merge793 (.A0(net64),
    .A1(net54),
    .A2(net50),
    .A3(net228),
    .S0(net101),
    .S1(net976),
    .X(net758));
 sky130_fd_sc_hd__clkbuf_1 merge794 (.A(net927),
    .X(net759));
 sky130_fd_sc_hd__mux4_1 merge795 (.A0(net278),
    .A1(clknet_1_1__leaf_net274),
    .A2(net983),
    .A3(net184),
    .S0(clknet_1_0__leaf_net291),
    .S1(clknet_1_1__leaf_net307),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_1 merge796 (.A(net822),
    .X(net761));
 sky130_fd_sc_hd__sedfxbp_1 merge797 (.CLK(clknet_4_1_0_clk),
    .D(net402),
    .DE(net404),
    .SCD(net539),
    .SCE(net417),
    .Q(net763),
    .Q_N(net762));
 sky130_fd_sc_hd__sdfbbn_1 merge798 (.CLK_N(clknet_4_15_0_clk),
    .D(clknet_1_1__leaf_net218),
    .RESET_B(net334),
    .SCD(net105),
    .SCE(net219),
    .SET_B(clknet_1_1__leaf_net971),
    .Q(net765),
    .Q_N(net764));
 sky130_fd_sc_hd__mux4_1 merge799 (.A0(net39),
    .A1(net284),
    .A2(net289),
    .A3(net288),
    .S0(net36),
    .S1(clknet_1_0__leaf_net841),
    .X(net766));
 sky130_fd_sc_hd__mux4_1 merge800 (.A0(net408),
    .A1(net265),
    .A2(net410),
    .A3(net954),
    .S0(clknet_1_1__leaf_net269),
    .S1(net262),
    .X(net767));
 sky130_fd_sc_hd__mux4_1 merge801 (.A0(net527),
    .A1(net417),
    .A2(net404),
    .A3(net530),
    .S0(net538),
    .S1(clknet_1_1__leaf_net537),
    .X(net768));
 sky130_fd_sc_hd__mux4_1 merge802 (.A0(clknet_1_1__leaf_net295),
    .A1(net245),
    .A2(net296),
    .A3(net276),
    .S0(net198),
    .S1(clknet_1_0__leaf_net843),
    .X(net769));
 sky130_fd_sc_hd__or4bb_1 merge803 (.A(net526),
    .B(net624),
    .C_N(net506),
    .D_N(net812),
    .X(net770));
 sky130_fd_sc_hd__mux4_1 merge804 (.A0(net55),
    .A1(net51),
    .A2(net53),
    .A3(net227),
    .S0(clknet_1_1__leaf_net815),
    .S1(net846),
    .X(net771));
 sky130_fd_sc_hd__mux4_1 merge805 (.A0(net275),
    .A1(net277),
    .A2(net287),
    .A3(net133),
    .S0(net156),
    .S1(net851),
    .X(net772));
 sky130_fd_sc_hd__or4bb_1 merge806 (.A(net627),
    .B(net621),
    .C_N(net526),
    .D_N(net1041),
    .X(net773));
 sky130_fd_sc_hd__mux4_1 merge807 (.A0(net630),
    .A1(net627),
    .A2(net998),
    .A3(net145),
    .S0(net21),
    .S1(clknet_1_0__leaf_net427),
    .X(net774));
 sky130_fd_sc_hd__sdfbbp_1 merge808 (.CLK(clknet_4_13_0_clk),
    .D(net53),
    .RESET_B(net15),
    .SCD(net46),
    .SCE(net1049),
    .SET_B(net57),
    .Q(net776),
    .Q_N(net775));
 sky130_fd_sc_hd__mux4_1 merge809 (.A0(net541),
    .A1(net404),
    .A2(net407),
    .A3(net76),
    .S0(clknet_1_0__leaf_net218),
    .S1(net319),
    .X(net777));
 sky130_fd_sc_hd__mux4_1 merge810 (.A0(net385),
    .A1(net381),
    .A2(net377),
    .A3(net625),
    .S0(net506),
    .S1(net796),
    .X(net778));
 sky130_fd_sc_hd__mux4_1 merge811 (.A0(net647),
    .A1(net506),
    .A2(net532),
    .A3(clknet_1_0__leaf_net537),
    .S0(net619),
    .S1(net998),
    .X(net779));
 sky130_fd_sc_hd__a2111o_1 merge812 (.A1(net522),
    .A2(net506),
    .B1(net1014),
    .C1(net1050),
    .D1(net1055),
    .X(net780));
 sky130_fd_sc_hd__dfrbp_1 merge813 (.CLK(clknet_4_13_0_clk),
    .D(net85),
    .RESET_B(net743),
    .Q(net782),
    .Q_N(net781));
 sky130_fd_sc_hd__dfrbp_1 merge814 (.CLK(clknet_4_6_0_clk),
    .D(net444),
    .RESET_B(net452),
    .Q(net784),
    .Q_N(net783));
 sky130_fd_sc_hd__dfrtn_1 merge815 (.CLK_N(clknet_4_15_0_clk),
    .D(net229),
    .RESET_B(net231),
    .Q(net785));
 sky130_fd_sc_hd__dfrtp_1 merge816 (.CLK(clknet_4_15_0_clk),
    .D(net360),
    .RESET_B(net361),
    .Q(net786));
 sky130_fd_sc_hd__dfrtp_1 merge817 (.CLK(clknet_4_2_0_clk),
    .D(net695),
    .RESET_B(net697),
    .Q(net787));
 sky130_fd_sc_hd__dfrtp_2 merge818 (.CLK(clknet_4_5_0_clk),
    .D(net160),
    .RESET_B(net173),
    .Q(net788));
 sky130_fd_sc_hd__dfsbp_1 merge819 (.CLK(clknet_4_14_0_clk),
    .D(net347),
    .SET_B(net353),
    .Q(net790),
    .Q_N(net789));
 sky130_fd_sc_hd__dfsbp_1 merge820 (.CLK(clknet_4_2_0_clk),
    .D(net665),
    .SET_B(net666),
    .Q(net792),
    .Q_N(net791));
 sky130_fd_sc_hd__dfstp_1 merge821 (.CLK(clknet_4_9_0_clk),
    .D(net465),
    .SET_B(net479),
    .Q(net793));
 sky130_fd_sc_hd__dfstp_1 merge822 (.CLK(clknet_4_4_0_clk),
    .D(net298),
    .SET_B(net752),
    .Q(net794));
 sky130_fd_sc_hd__dfstp_1 merge823 (.CLK(clknet_4_1_0_clk),
    .D(net396),
    .SET_B(net392),
    .Q(net795));
 sky130_fd_sc_hd__dlrbn_1 merge824 (.D(net648),
    .GATE_N(clknet_4_0_0_clk),
    .RESET_B(net652),
    .Q(net797),
    .Q_N(net796));
 sky130_fd_sc_hd__dlrbn_1 merge825 (.D(net568),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net570),
    .Q(net799),
    .Q_N(net798));
 sky130_fd_sc_hd__dlrbp_1 merge826 (.D(net595),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net597),
    .Q(net801),
    .Q_N(net800));
 sky130_fd_sc_hd__dlrbp_1 merge827 (.D(net729),
    .GATE(clknet_4_0_0_clk),
    .RESET_B(net770),
    .Q(net803),
    .Q_N(net802));
 sky130_fd_sc_hd__dlrtn_2 merge828 (.D(net727),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net756),
    .Q(net804));
 sky130_fd_sc_hd__dlrtn_1 merge829 (.D(net504),
    .GATE_N(clknet_4_11_0_clk),
    .RESET_B(net498),
    .Q(net805));
 sky130_fd_sc_hd__dlrtn_1 merge830 (.D(net710),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net713),
    .Q(net806));
 sky130_fd_sc_hd__dlrtp_2 merge831 (.D(net734),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net92),
    .Q(net807));
 sky130_fd_sc_hd__dlrtp_1 merge832 (.D(net207),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net745),
    .Q(net808));
 sky130_fd_sc_hd__dlrtp_1 merge833 (.D(net412),
    .GATE(clknet_4_1_0_clk),
    .Q(net413));
 sky130_fd_sc_hd__edfxbp_1 merge834 (.CLK(clknet_4_3_0_clk),
    .D(net576),
    .DE(net580),
    .Q(net811),
    .Q_N(net810));
 sky130_fd_sc_hd__edfxtp_1 merge835 (.CLK(clknet_4_0_0_clk),
    .D(net525),
    .DE(net523),
    .Q(net812));
 sky130_fd_sc_hd__sdlclkp_1 merge836 (.CLK(clknet_4_13_0_clk),
    .GATE(net179),
    .SCE(net188),
    .GCLK(net813));
 sky130_fd_sc_hd__sdlclkp_2 merge837 (.CLK(clknet_4_4_0_clk),
    .GATE(net279),
    .SCE(net746),
    .GCLK(net814));
 sky130_fd_sc_hd__sdlclkp_4 merge838 (.CLK(clknet_4_5_0_clk),
    .GATE(net152),
    .SCE(net144),
    .GCLK(net815));
 sky130_fd_sc_hd__dfrbp_1 merge839 (.CLK(clknet_4_1_0_clk),
    .D(net545),
    .RESET_B(net744),
    .Q(net817),
    .Q_N(net816));
 sky130_fd_sc_hd__dfrbp_1 merge840 (.CLK(clknet_4_12_0_clk),
    .D(net324),
    .RESET_B(net325),
    .Q(net819),
    .Q_N(net818));
 sky130_fd_sc_hd__dfrtn_1 merge841 (.CLK_N(clknet_4_6_0_clk),
    .D(net434),
    .RESET_B(net428),
    .Q(net820));
 sky130_fd_sc_hd__dfrtp_1 merge842 (.CLK(clknet_4_11_0_clk),
    .D(net592),
    .RESET_B(net500),
    .Q(net821));
 sky130_fd_sc_hd__dfrtp_4 merge843 (.CLK(clknet_4_0_0_clk),
    .D(net777),
    .RESET_B(net780),
    .Q(net822));
 sky130_fd_sc_hd__dfrtp_1 merge844 (.CLK(clknet_4_4_0_clk),
    .D(net416),
    .RESET_B(net437),
    .Q(net823));
 sky130_fd_sc_hd__dfsbp_1 merge845 (.CLK(clknet_4_8_0_clk),
    .D(net700),
    .SET_B(net722),
    .Q(net825),
    .Q_N(net824));
 sky130_fd_sc_hd__dfsbp_1 merge846 (.CLK(clknet_4_2_0_clk),
    .D(net684),
    .SET_B(net705),
    .Q(net827),
    .Q_N(net826));
 sky130_fd_sc_hd__dfstp_1 merge847 (.CLK(clknet_4_10_0_clk),
    .D(net702),
    .SET_B(net499),
    .Q(net828));
 sky130_fd_sc_hd__dfstp_1 merge848 (.CLK(clknet_4_11_0_clk),
    .D(net599),
    .SET_B(net600),
    .Q(net972));
 sky130_fd_sc_hd__dfstp_1 merge849 (.CLK(clknet_4_11_0_clk),
    .D(net611),
    .SET_B(net457),
    .Q(net829));
 sky130_fd_sc_hd__dlrbn_1 merge850 (.D(net742),
    .GATE_N(clknet_4_0_0_clk),
    .RESET_B(net773),
    .Q(net831),
    .Q_N(net830));
 sky130_fd_sc_hd__dlrbn_1 merge851 (.D(net149),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net148),
    .Q(net833),
    .Q_N(net832));
 sky130_fd_sc_hd__dfxbp_1 s852 (.CLK(clknet_4_7_0_clk),
    .D(net38),
    .Q(net835),
    .Q_N(net834));
 sky130_fd_sc_hd__dfxbp_1 s853 (.CLK(clknet_4_13_0_clk),
    .D(net60),
    .Q(net837),
    .Q_N(net836));
 sky130_fd_sc_hd__dfxtp_1 s854 (.CLK(clknet_4_13_0_clk),
    .D(net62),
    .Q(net838));
 sky130_fd_sc_hd__dfxtp_1 s855 (.CLK(clknet_4_15_0_clk),
    .D(net86),
    .Q(net839));
 sky130_fd_sc_hd__dfxtp_1 s856 (.CLK(clknet_4_5_0_clk),
    .D(net171),
    .Q(net840));
 sky130_fd_sc_hd__dlclkp_1 s857 (.CLK(clknet_4_13_0_clk),
    .GATE(net189),
    .GCLK(net841));
 sky130_fd_sc_hd__dlclkp_2 s858 (.CLK(clknet_4_12_0_clk),
    .GATE(net195),
    .GCLK(net842));
 sky130_fd_sc_hd__dlclkp_4 s859 (.CLK(clknet_4_12_0_clk),
    .GATE(net196),
    .GCLK(net843));
 sky130_fd_sc_hd__dlxbn_1 s860 (.D(net224),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net845),
    .Q_N(net844));
 sky130_fd_sc_hd__dlxbn_1 s861 (.D(net233),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net847),
    .Q_N(net846));
 sky130_fd_sc_hd__dlxbp_1 s862 (.D(net237),
    .GATE(clknet_4_15_0_clk),
    .Q(net849),
    .Q_N(net848));
 sky130_fd_sc_hd__dlxtn_1 s863 (.D(net238),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net850));
 sky130_fd_sc_hd__dlxtn_1 s864 (.D(net272),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net851));
 sky130_fd_sc_hd__dlxtn_4 s865 (.D(net299),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net852));
 sky130_fd_sc_hd__dlxtp_1 s866 (.D(net300),
    .GATE(clknet_4_6_0_clk),
    .Q(net853));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s867 (.D(net309),
    .SLEEP_B(clknet_4_12_0_clk),
    .Q(net854));
 sky130_fd_sc_hd__dfxbp_1 s868 (.CLK(clknet_4_12_0_clk),
    .D(net312),
    .Q(net856),
    .Q_N(net855));
 sky130_fd_sc_hd__dfxbp_1 s869 (.CLK(clknet_4_14_0_clk),
    .D(net326),
    .Q(net857));
 sky130_fd_sc_hd__dfxtp_1 s870 (.CLK(clknet_4_14_0_clk),
    .D(net349),
    .Q(net858));
 sky130_fd_sc_hd__dfxtp_1 s871 (.CLK(clknet_4_15_0_clk),
    .D(net363),
    .Q(net859));
 sky130_fd_sc_hd__dfxtp_1 s872 (.CLK(clknet_4_14_0_clk),
    .D(net369),
    .Q(net860));
 sky130_fd_sc_hd__dlclkp_1 s873 (.CLK(clknet_4_14_0_clk),
    .GATE(net370),
    .GCLK(net861));
 sky130_fd_sc_hd__dlclkp_2 s874 (.CLK(clknet_4_11_0_clk),
    .GATE(net371),
    .GCLK(net862));
 sky130_fd_sc_hd__dlclkp_4 s875 (.CLK(clknet_4_14_0_clk),
    .GATE(net372),
    .GCLK(net863));
 sky130_fd_sc_hd__dlxbn_1 s876 (.D(net414),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net865),
    .Q_N(net864));
 sky130_fd_sc_hd__dlxbn_1 s877 (.D(net418),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net867),
    .Q_N(net866));
 sky130_fd_sc_hd__dlxbp_1 s878 (.D(net433),
    .GATE(clknet_4_3_0_clk),
    .Q(net869),
    .Q_N(net868));
 sky130_fd_sc_hd__dlxtn_2 s879 (.D(net436),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net870));
 sky130_fd_sc_hd__dlxtn_1 s880 (.D(net454),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net871));
 sky130_fd_sc_hd__dlxtn_1 s881 (.D(net461),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net872));
 sky130_fd_sc_hd__dlxtp_1 s882 (.D(net462),
    .GATE(clknet_4_9_0_clk),
    .Q(net873));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s883 (.D(net472),
    .SLEEP_B(clknet_4_11_0_clk),
    .Q(net874));
 sky130_fd_sc_hd__dfxbp_1 s884 (.CLK(clknet_4_11_0_clk),
    .D(net476),
    .Q(net876),
    .Q_N(net875));
 sky130_fd_sc_hd__dfxbp_1 s885 (.CLK(clknet_4_14_0_clk),
    .D(net484),
    .Q(net878),
    .Q_N(net877));
 sky130_fd_sc_hd__dfxtp_2 s886 (.CLK(clknet_4_11_0_clk),
    .D(net496),
    .Q(net879));
 sky130_fd_sc_hd__dfxtp_2 s887 (.CLK(clknet_4_3_0_clk),
    .D(net564),
    .Q(net880));
 sky130_fd_sc_hd__dfxtp_2 s888 (.CLK(clknet_4_2_0_clk),
    .D(net571),
    .Q(net881));
 sky130_fd_sc_hd__dlclkp_1 s889 (.CLK(clknet_4_3_0_clk),
    .GATE(net572),
    .GCLK(net882));
 sky130_fd_sc_hd__dlclkp_2 s890 (.CLK(clknet_4_3_0_clk),
    .GATE(net581),
    .GCLK(net963));
 sky130_fd_sc_hd__dlclkp_4 s891 (.CLK(clknet_4_3_0_clk),
    .GATE(net582),
    .GCLK(net883));
 sky130_fd_sc_hd__dlxbn_1 s892 (.D(net586),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net885),
    .Q_N(net884));
 sky130_fd_sc_hd__dlxbn_1 s893 (.D(net588),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net887),
    .Q_N(net886));
 sky130_fd_sc_hd__dlxbp_1 s894 (.D(net590),
    .GATE(clknet_4_8_0_clk),
    .Q(net889),
    .Q_N(net888));
 sky130_fd_sc_hd__dlxtn_2 s895 (.D(net591),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net890));
 sky130_fd_sc_hd__dlxtn_1 s896 (.D(net593),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net891));
 sky130_fd_sc_hd__dlxtn_1 s897 (.D(net598),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net892));
 sky130_fd_sc_hd__dlxtp_1 s898 (.D(net613),
    .GATE(clknet_4_10_0_clk),
    .Q(net893));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s899 (.D(net651),
    .SLEEP_B(clknet_4_0_0_clk),
    .Q(net894));
 sky130_fd_sc_hd__dfxbp_1 s900 (.CLK(clknet_4_8_0_clk),
    .D(net682),
    .Q(net896),
    .Q_N(net895));
 sky130_fd_sc_hd__dfxbp_1 s901 (.CLK(clknet_4_2_0_clk),
    .D(net683),
    .Q(net898),
    .Q_N(net897));
 sky130_fd_sc_hd__dfxtp_1 s902 (.CLK(clknet_4_2_0_clk),
    .D(net686),
    .Q(net899));
 sky130_fd_sc_hd__dfxtp_1 s903 (.CLK(clknet_4_8_0_clk),
    .D(net694),
    .Q(net900));
 sky130_fd_sc_hd__dfxtp_2 s904 (.CLK(clknet_4_2_0_clk),
    .D(net701),
    .Q(net901));
 sky130_fd_sc_hd__dlclkp_1 s905 (.CLK(clknet_4_8_0_clk),
    .GATE(net703),
    .GCLK(net902));
 sky130_fd_sc_hd__dlclkp_2 s906 (.CLK(clknet_4_8_0_clk),
    .GATE(net704),
    .GCLK(net903));
 sky130_fd_sc_hd__dlclkp_4 s907 (.CLK(clknet_4_8_0_clk),
    .GATE(net706),
    .GCLK(net904));
 sky130_fd_sc_hd__dlxbn_1 s908 (.D(net707),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net906),
    .Q_N(net905));
 sky130_fd_sc_hd__dlxbn_1 s909 (.D(net717),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net907));
 sky130_fd_sc_hd__dlxbp_1 s910 (.D(net718),
    .GATE(clknet_4_8_0_clk),
    .Q(net909),
    .Q_N(net908));
 sky130_fd_sc_hd__dlxtn_1 s911 (.D(net720),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net910));
 sky130_fd_sc_hd__dlxtn_1 s912 (.D(net725),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net911));
 sky130_fd_sc_hd__dlxtn_1 s913 (.D(net726),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net912));
 sky130_fd_sc_hd__dlxtp_1 s914 (.D(net728),
    .GATE(clknet_4_0_0_clk),
    .Q(net913));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s915 (.D(net733),
    .SLEEP_B(clknet_4_13_0_clk),
    .Q(net914));
 sky130_fd_sc_hd__dfxbp_1 s916 (.CLK(clknet_4_6_0_clk),
    .D(net740),
    .Q(net916),
    .Q_N(net915));
 sky130_fd_sc_hd__dfxbp_1 s917 (.CLK(clknet_4_2_0_clk),
    .D(net753),
    .Q(net918),
    .Q_N(net917));
 sky130_fd_sc_hd__dfxtp_1 s918 (.CLK(clknet_4_4_0_clk),
    .D(net755),
    .Q(net919));
 sky130_fd_sc_hd__dfxtp_1 s919 (.CLK(clknet_4_13_0_clk),
    .D(net757),
    .Q(net920));
 sky130_fd_sc_hd__dfxtp_1 s920 (.CLK(clknet_4_15_0_clk),
    .D(net758),
    .Q(net921));
 sky130_fd_sc_hd__dlclkp_1 s921 (.CLK(clknet_4_7_0_clk),
    .GATE(net760),
    .GCLK(net922));
 sky130_fd_sc_hd__dlclkp_2 s922 (.CLK(clknet_4_7_0_clk),
    .GATE(net766),
    .GCLK(net923));
 sky130_fd_sc_hd__dlclkp_4 s923 (.CLK(clknet_4_4_0_clk),
    .GATE(net767),
    .GCLK(net924));
 sky130_fd_sc_hd__dlxbn_1 s924 (.D(net768),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net926),
    .Q_N(net925));
 sky130_fd_sc_hd__dlxbn_1 s925 (.D(net769),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net928),
    .Q_N(net927));
 sky130_fd_sc_hd__dlxbp_1 s926 (.D(net771),
    .GATE(clknet_4_13_0_clk),
    .Q(net930),
    .Q_N(net929));
 sky130_fd_sc_hd__dlxtn_1 s927 (.D(net772),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net931));
 sky130_fd_sc_hd__dlxtn_1 s928 (.D(net774),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net932));
 sky130_fd_sc_hd__dlxtn_1 s929 (.D(net778),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net933));
 sky130_fd_sc_hd__dlxtp_1 s930 (.D(net779),
    .GATE(clknet_4_0_0_clk),
    .Q(net934));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(in0),
    .X(net738));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(in1),
    .X(net935));
 sky130_fd_sc_hd__buf_4 input3 (.A(in10),
    .X(net936));
 sky130_fd_sc_hd__buf_2 input4 (.A(in11),
    .X(net937));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(in12),
    .X(net938));
 sky130_fd_sc_hd__buf_2 input6 (.A(in13),
    .X(net939));
 sky130_fd_sc_hd__buf_1 input7 (.A(in14),
    .X(net940));
 sky130_fd_sc_hd__buf_2 input8 (.A(in15),
    .X(net941));
 sky130_fd_sc_hd__buf_4 input9 (.A(in16),
    .X(net942));
 sky130_fd_sc_hd__buf_2 input10 (.A(in17),
    .X(net943));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(in18),
    .X(net944));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(in19),
    .X(net945));
 sky130_fd_sc_hd__buf_1 input13 (.A(in2),
    .X(net946));
 sky130_fd_sc_hd__buf_1 input14 (.A(in20),
    .X(net947));
 sky130_fd_sc_hd__buf_1 input15 (.A(in21),
    .X(net948));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(in22),
    .X(net949));
 sky130_fd_sc_hd__buf_4 input17 (.A(in23),
    .X(net950));
 sky130_fd_sc_hd__buf_2 input18 (.A(in24),
    .X(net951));
 sky130_fd_sc_hd__buf_1 input19 (.A(in3),
    .X(net952));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(in4),
    .X(net953));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(in5),
    .X(net954));
 sky130_fd_sc_hd__buf_2 input22 (.A(in6),
    .X(net955));
 sky130_fd_sc_hd__buf_2 input23 (.A(in7),
    .X(net956));
 sky130_fd_sc_hd__buf_4 input24 (.A(in8),
    .X(net957));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(in9),
    .X(net958));
 sky130_fd_sc_hd__buf_2 output26 (.A(net959),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output27 (.A(net960),
    .X(out1));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(clknet_1_1__leaf_net961),
    .X(out10));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(clknet_1_1__leaf_net962),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(clknet_1_0__leaf_net963),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output31 (.A(net989),
    .X(out13));
 sky130_fd_sc_hd__clkbuf_1 output32 (.A(clknet_1_0__leaf_net965),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output33 (.A(net966),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output34 (.A(net967),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output35 (.A(net992),
    .X(out17));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(clknet_1_1__leaf_net969),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output37 (.A(net970),
    .X(out19));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(clknet_1_0__leaf_net971),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output39 (.A(net972),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output40 (.A(net973),
    .X(out21));
 sky130_fd_sc_hd__clkbuf_1 output41 (.A(net974),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output42 (.A(net987),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output43 (.A(net976),
    .X(out24));
 sky130_fd_sc_hd__clkbuf_1 output44 (.A(clknet_1_1__leaf_net977),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output45 (.A(net978),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output46 (.A(net979),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output47 (.A(net980),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output48 (.A(net981),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_1 output49 (.A(clknet_1_0__leaf_net982),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output50 (.A(net983),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_4 fanout51 (.A(net185),
    .X(net984));
 sky130_fd_sc_hd__buf_2 fanout52 (.A(net680),
    .X(net985));
 sky130_fd_sc_hd__buf_4 fanout53 (.A(net975),
    .X(net986));
 sky130_fd_sc_hd__clkbuf_2 fanout54 (.A(net975),
    .X(net987));
 sky130_fd_sc_hd__buf_2 fanout55 (.A(net512),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_4 fanout56 (.A(net964),
    .X(net989));
 sky130_fd_sc_hd__clkbuf_2 fanout57 (.A(net964),
    .X(net990));
 sky130_fd_sc_hd__clkbuf_4 fanout58 (.A(net405),
    .X(net991));
 sky130_fd_sc_hd__buf_4 fanout59 (.A(net968),
    .X(net992));
 sky130_fd_sc_hd__clkbuf_4 fanout60 (.A(net264),
    .X(net993));
 sky130_fd_sc_hd__buf_4 fanout61 (.A(net259),
    .X(net994));
 sky130_fd_sc_hd__clkbuf_4 fanout62 (.A(net165),
    .X(net995));
 sky130_fd_sc_hd__clkbuf_4 fanout63 (.A(net77),
    .X(net996));
 sky130_fd_sc_hd__clkbuf_4 fanout64 (.A(net115),
    .X(net997));
 sky130_fd_sc_hd__buf_2 fanout65 (.A(net999),
    .X(net998));
 sky130_fd_sc_hd__clkbuf_2 fanout66 (.A(net629),
    .X(net999));
 sky130_fd_sc_hd__clkbuf_4 fanout67 (.A(net552),
    .X(net1000));
 sky130_fd_sc_hd__buf_2 fanout68 (.A(net223),
    .X(net1001));
 sky130_fd_sc_hd__buf_4 fanout69 (.A(net873),
    .X(net1002));
 sky130_fd_sc_hd__clkbuf_4 fanout70 (.A(net868),
    .X(net1003));
 sky130_fd_sc_hd__buf_4 fanout71 (.A(net869),
    .X(net1004));
 sky130_fd_sc_hd__clkbuf_2 fanout72 (.A(net869),
    .X(net1005));
 sky130_fd_sc_hd__clkbuf_4 fanout73 (.A(net981),
    .X(net1006));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net924 (.A(net924),
    .X(clknet_0_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net924 (.A(clknet_0_net924),
    .X(clknet_1_0__leaf_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net924 (.A(clknet_0_net924),
    .X(clknet_1_1__leaf_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net415 (.A(net415),
    .X(clknet_0_net415));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net415 (.A(clknet_0_net415),
    .X(clknet_1_0__leaf_net415));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net415 (.A(clknet_0_net415),
    .X(clknet_1_1__leaf_net415));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net555 (.A(net555),
    .X(clknet_0_net555));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net555 (.A(clknet_0_net555),
    .X(clknet_1_0__leaf_net555));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net555 (.A(clknet_0_net555),
    .X(clknet_1_1__leaf_net555));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net883 (.A(net883),
    .X(clknet_0_net883));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net883 (.A(clknet_0_net883),
    .X(clknet_1_0__leaf_net883));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net883 (.A(clknet_0_net883),
    .X(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net589 (.A(net589),
    .X(clknet_0_net589));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net589 (.A(clknet_0_net589),
    .X(clknet_1_0__leaf_net589));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net589 (.A(clknet_0_net589),
    .X(clknet_1_1__leaf_net589));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net587 (.A(net587),
    .X(clknet_0_net587));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net587 (.A(clknet_0_net587),
    .X(clknet_1_0__leaf_net587));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net587 (.A(clknet_0_net587),
    .X(clknet_1_1__leaf_net587));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net584 (.A(net584),
    .X(clknet_0_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net584 (.A(clknet_0_net584),
    .X(clknet_1_0__leaf_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net584 (.A(clknet_0_net584),
    .X(clknet_1_1__leaf_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net961 (.A(net961),
    .X(clknet_0_net961));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net961 (.A(clknet_0_net961),
    .X(clknet_1_0__leaf_net961));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net961 (.A(clknet_0_net961),
    .X(clknet_1_1__leaf_net961));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net583 (.A(net583),
    .X(clknet_0_net583));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net583 (.A(clknet_0_net583),
    .X(clknet_1_0__leaf_net583));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net583 (.A(clknet_0_net583),
    .X(clknet_1_1__leaf_net583));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net982 (.A(net982),
    .X(clknet_0_net982));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net982 (.A(clknet_0_net982),
    .X(clknet_1_0__leaf_net982));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net982 (.A(clknet_0_net982),
    .X(clknet_1_1__leaf_net982));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net273 (.A(net273),
    .X(clknet_0_net273));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net273 (.A(clknet_0_net273),
    .X(clknet_1_0__leaf_net273));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net273 (.A(clknet_0_net273),
    .X(clknet_1_1__leaf_net273));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net281 (.A(net281),
    .X(clknet_0_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net281 (.A(clknet_0_net281),
    .X(clknet_1_0__leaf_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net281 (.A(clknet_0_net281),
    .X(clknet_1_1__leaf_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net411 (.A(net411),
    .X(clknet_0_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net411 (.A(clknet_0_net411),
    .X(clknet_1_0__leaf_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net411 (.A(clknet_0_net411),
    .X(clknet_1_1__leaf_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net553 (.A(net553),
    .X(clknet_0_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net553 (.A(clknet_0_net553),
    .X(clknet_1_0__leaf_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net553 (.A(clknet_0_net553),
    .X(clknet_1_1__leaf_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net274 (.A(net274),
    .X(clknet_0_net274));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net274 (.A(clknet_0_net274),
    .X(clknet_1_0__leaf_net274));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net274 (.A(clknet_0_net274),
    .X(clknet_1_1__leaf_net274));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net922 (.A(net922),
    .X(clknet_0_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net922 (.A(clknet_0_net922),
    .X(clknet_1_0__leaf_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net922 (.A(clknet_0_net922),
    .X(clknet_1_1__leaf_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net327 (.A(net327),
    .X(clknet_0_net327));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net327 (.A(clknet_0_net327),
    .X(clknet_1_0__leaf_net327));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net327 (.A(clknet_0_net327),
    .X(clknet_1_1__leaf_net327));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net491 (.A(net491),
    .X(clknet_0_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net491 (.A(clknet_0_net491),
    .X(clknet_1_0__leaf_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net491 (.A(clknet_0_net491),
    .X(clknet_1_1__leaf_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net497 (.A(net497),
    .X(clknet_0_net497));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net497 (.A(clknet_0_net497),
    .X(clknet_1_0__leaf_net497));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net497 (.A(clknet_0_net497),
    .X(clknet_1_1__leaf_net497));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net485 (.A(net485),
    .X(clknet_0_net485));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net485 (.A(clknet_0_net485),
    .X(clknet_1_0__leaf_net485));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net485 (.A(clknet_0_net485),
    .X(clknet_1_1__leaf_net485));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net453 (.A(net453),
    .X(clknet_0_net453));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net453 (.A(clknet_0_net453),
    .X(clknet_1_0__leaf_net453));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net453 (.A(clknet_0_net453),
    .X(clknet_1_1__leaf_net453));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net969 (.A(net969),
    .X(clknet_0_net969));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net969 (.A(clknet_0_net969),
    .X(clknet_1_0__leaf_net969));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net969 (.A(clknet_0_net969),
    .X(clknet_1_1__leaf_net969));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net280 (.A(net280),
    .X(clknet_0_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net280 (.A(clknet_0_net280),
    .X(clknet_1_0__leaf_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net280 (.A(clknet_0_net280),
    .X(clknet_1_1__leaf_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net291 (.A(net291),
    .X(clknet_0_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net291 (.A(clknet_0_net291),
    .X(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net291 (.A(clknet_0_net291),
    .X(clknet_1_1__leaf_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net314 (.A(net314),
    .X(clknet_0_net314));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net314 (.A(net1010),
    .X(clknet_1_0__leaf_net314));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net314 (.A(clknet_0_net314),
    .X(clknet_1_1__leaf_net314));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net882 (.A(net882),
    .X(clknet_0_net882));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net882 (.A(clknet_0_net882),
    .X(clknet_1_0__leaf_net882));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net882 (.A(clknet_0_net882),
    .X(clknet_1_1__leaf_net882));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net328 (.A(net328),
    .X(clknet_0_net328));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net328 (.A(net1011),
    .X(clknet_1_0__leaf_net328));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net328 (.A(clknet_0_net328),
    .X(clknet_1_1__leaf_net328));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net473 (.A(net473),
    .X(clknet_0_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net473 (.A(clknet_0_net473),
    .X(clknet_1_0__leaf_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net473 (.A(clknet_0_net473),
    .X(clknet_1_1__leaf_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net456 (.A(net456),
    .X(clknet_0_net456));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net456 (.A(clknet_0_net456),
    .X(clknet_1_0__leaf_net456));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net456 (.A(clknet_0_net456),
    .X(clknet_1_1__leaf_net456));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net923 (.A(net923),
    .X(clknet_0_net923));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net923 (.A(clknet_0_net923),
    .X(clknet_1_0__leaf_net923));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net923 (.A(clknet_0_net923),
    .X(clknet_1_1__leaf_net923));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net307 (.A(net307),
    .X(clknet_0_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net307 (.A(clknet_0_net307),
    .X(clknet_1_0__leaf_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net307 (.A(clknet_0_net307),
    .X(clknet_1_1__leaf_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net451 (.A(net451),
    .X(clknet_0_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net451 (.A(clknet_0_net451),
    .X(clknet_1_0__leaf_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net451 (.A(clknet_0_net451),
    .X(clknet_1_1__leaf_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net450 (.A(net450),
    .X(clknet_0_net450));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net450 (.A(clknet_0_net450),
    .X(clknet_1_0__leaf_net450));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net450 (.A(clknet_0_net450),
    .X(clknet_1_1__leaf_net450));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net963 (.A(net963),
    .X(clknet_0_net963));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net963 (.A(clknet_0_net963),
    .X(clknet_1_0__leaf_net963));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net963 (.A(clknet_0_net963),
    .X(clknet_1_1__leaf_net963));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net460 (.A(net460),
    .X(clknet_0_net460));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net460 (.A(clknet_0_net460),
    .X(clknet_1_0__leaf_net460));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net460 (.A(clknet_0_net460),
    .X(clknet_1_1__leaf_net460));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net441 (.A(net441),
    .X(clknet_0_net441));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net441 (.A(clknet_0_net441),
    .X(clknet_1_0__leaf_net441));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net441 (.A(clknet_0_net441),
    .X(clknet_1_1__leaf_net441));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net698 (.A(net698),
    .X(clknet_0_net698));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net698 (.A(clknet_0_net698),
    .X(clknet_1_0__leaf_net698));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net698 (.A(clknet_0_net698),
    .X(clknet_1_1__leaf_net698));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net904 (.A(net904),
    .X(clknet_0_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net904 (.A(clknet_0_net904),
    .X(clknet_1_0__leaf_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net904 (.A(clknet_0_net904),
    .X(clknet_1_1__leaf_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net708 (.A(net708),
    .X(clknet_0_net708));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net708 (.A(clknet_0_net708),
    .X(clknet_1_0__leaf_net708));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net708 (.A(clknet_0_net708),
    .X(clknet_1_1__leaf_net708));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net316 (.A(net316),
    .X(clknet_0_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net316 (.A(clknet_0_net316),
    .X(clknet_1_0__leaf_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net316 (.A(clknet_0_net316),
    .X(clknet_1_1__leaf_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net295 (.A(net295),
    .X(clknet_0_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net295 (.A(clknet_0_net295),
    .X(clknet_1_0__leaf_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net295 (.A(clknet_0_net295),
    .X(clknet_1_1__leaf_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net863 (.A(net863),
    .X(clknet_0_net863));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net863 (.A(clknet_0_net863),
    .X(clknet_1_0__leaf_net863));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net863 (.A(clknet_0_net863),
    .X(clknet_1_1__leaf_net863));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net862 (.A(net862),
    .X(clknet_0_net862));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net862 (.A(clknet_0_net862),
    .X(clknet_1_0__leaf_net862));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net862 (.A(clknet_0_net862),
    .X(clknet_1_1__leaf_net862));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net843 (.A(net843),
    .X(clknet_0_net843));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net843 (.A(clknet_0_net843),
    .X(clknet_1_0__leaf_net843));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net843 (.A(clknet_0_net843),
    .X(clknet_1_1__leaf_net843));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net310 (.A(net310),
    .X(clknet_0_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net310 (.A(clknet_0_net310),
    .X(clknet_1_0__leaf_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net310 (.A(clknet_0_net310),
    .X(clknet_1_1__leaf_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net197 (.A(net197),
    .X(clknet_0_net197));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net197 (.A(clknet_0_net197),
    .X(clknet_1_0__leaf_net197));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net197 (.A(clknet_0_net197),
    .X(clknet_1_1__leaf_net197));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net217 (.A(net217),
    .X(clknet_0_net217));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net217 (.A(clknet_0_net217),
    .X(clknet_1_0__leaf_net217));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net217 (.A(clknet_0_net217),
    .X(clknet_1_1__leaf_net217));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net348 (.A(net348),
    .X(clknet_0_net348));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net348 (.A(clknet_0_net348),
    .X(clknet_1_0__leaf_net348));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net348 (.A(clknet_0_net348),
    .X(clknet_1_1__leaf_net348));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net218 (.A(net218),
    .X(clknet_0_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net218 (.A(clknet_0_net218),
    .X(clknet_1_0__leaf_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net218 (.A(clknet_0_net218),
    .X(clknet_1_1__leaf_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net212 (.A(net212),
    .X(clknet_0_net212));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net212 (.A(clknet_0_net212),
    .X(clknet_1_0__leaf_net212));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net212 (.A(clknet_0_net212),
    .X(clknet_1_1__leaf_net212));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net962 (.A(net962),
    .X(clknet_0_net962));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net962 (.A(clknet_0_net962),
    .X(clknet_1_0__leaf_net962));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net962 (.A(clknet_0_net962),
    .X(clknet_1_1__leaf_net962));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net345 (.A(net345),
    .X(clknet_0_net345));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net345 (.A(clknet_0_net345),
    .X(clknet_1_0__leaf_net345));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net345 (.A(clknet_0_net345),
    .X(clknet_1_1__leaf_net345));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net842 (.A(net842),
    .X(clknet_0_net842));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net842 (.A(clknet_0_net842),
    .X(clknet_1_0__leaf_net842));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net842 (.A(clknet_0_net842),
    .X(clknet_1_1__leaf_net842));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net965 (.A(net965),
    .X(clknet_0_net965));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net965 (.A(clknet_0_net965),
    .X(clknet_1_0__leaf_net965));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net965 (.A(clknet_0_net965),
    .X(clknet_1_1__leaf_net965));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net841 (.A(net841),
    .X(clknet_0_net841));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net841 (.A(clknet_0_net841),
    .X(clknet_1_0__leaf_net841));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net841 (.A(clknet_0_net841),
    .X(clknet_1_1__leaf_net841));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net192 (.A(net192),
    .X(clknet_0_net192));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net192 (.A(clknet_0_net192),
    .X(clknet_1_0__leaf_net192));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net192 (.A(clknet_0_net192),
    .X(clknet_1_1__leaf_net192));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net815 (.A(net815),
    .X(clknet_0_net815));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net815 (.A(clknet_0_net815),
    .X(clknet_1_0__leaf_net815));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net815 (.A(clknet_0_net815),
    .X(clknet_1_1__leaf_net815));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net202 (.A(net202),
    .X(clknet_0_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net202 (.A(clknet_0_net202),
    .X(clknet_1_0__leaf_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net202 (.A(clknet_0_net202),
    .X(clknet_1_1__leaf_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net203 (.A(net203),
    .X(clknet_0_net203));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net203 (.A(clknet_0_net203),
    .X(clknet_1_0__leaf_net203));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net203 (.A(clknet_0_net203),
    .X(clknet_1_1__leaf_net203));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net971 (.A(net971),
    .X(clknet_0_net971));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net971 (.A(clknet_0_net971),
    .X(clknet_1_0__leaf_net971));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net971 (.A(clknet_0_net971),
    .X(clknet_1_1__leaf_net971));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net172 (.A(net172),
    .X(clknet_0_net172));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net172 (.A(clknet_0_net172),
    .X(clknet_1_0__leaf_net172));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net172 (.A(clknet_0_net172),
    .X(clknet_1_1__leaf_net172));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net294 (.A(net294),
    .X(clknet_0_net294));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net294 (.A(clknet_0_net294),
    .X(clknet_1_0__leaf_net294));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net294 (.A(clknet_0_net294),
    .X(clknet_1_1__leaf_net294));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net427 (.A(net427),
    .X(clknet_0_net427));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net427 (.A(clknet_0_net427),
    .X(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net427 (.A(clknet_0_net427),
    .X(clknet_1_1__leaf_net427));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net315 (.A(net315),
    .X(clknet_0_net315));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net315 (.A(clknet_0_net315),
    .X(clknet_1_0__leaf_net315));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net315 (.A(clknet_0_net315),
    .X(clknet_1_1__leaf_net315));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net977 (.A(net977),
    .X(clknet_0_net977));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net977 (.A(clknet_0_net977),
    .X(clknet_1_0__leaf_net977));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net977 (.A(clknet_0_net977),
    .X(clknet_1_1__leaf_net977));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net814 (.A(net814),
    .X(clknet_0_net814));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net814 (.A(clknet_0_net814),
    .X(clknet_1_0__leaf_net814));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net814 (.A(clknet_0_net814),
    .X(clknet_1_1__leaf_net814));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net269 (.A(net269),
    .X(clknet_0_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net269 (.A(clknet_0_net269),
    .X(clknet_1_0__leaf_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net269 (.A(clknet_0_net269),
    .X(clknet_1_1__leaf_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net537 (.A(net537),
    .X(clknet_0_net537));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net537 (.A(clknet_0_net537),
    .X(clknet_1_0__leaf_net537));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net537 (.A(clknet_0_net537),
    .X(clknet_1_1__leaf_net537));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net263 (.A(net263),
    .X(clknet_0_net263));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net263 (.A(clknet_0_net263),
    .X(clknet_1_0__leaf_net263));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net263 (.A(clknet_0_net263),
    .X(clknet_1_1__leaf_net263));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net813 (.A(net813),
    .X(clknet_0_net813));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net813 (.A(clknet_0_net813),
    .X(clknet_1_0__leaf_net813));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net813 (.A(clknet_0_net813),
    .X(clknet_1_1__leaf_net813));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net59),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net1007),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net1008),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(clknet_0_net314),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(clknet_0_net328),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net879),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net853),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net644),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net900),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net840),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net838),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net823),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net236),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net391),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net455),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net609),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net387),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net795),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net921),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net532),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net150),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net918),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net543),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net881),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net635),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net606),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net801),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net898),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net959),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net786),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net161),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net352),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net821),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net852),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net620),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net788),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net920),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net837),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net615),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net892),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net894),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net791),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net58),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net619),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net835),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net563),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net788),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net880),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net643),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net643),
    .X(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c54_B (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c35_B (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A0 (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c25_X (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S0 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_S0 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_A2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c28_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_X (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A0 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_S1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_C (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c35_X (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A3 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_S0 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A0 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_S1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_C_N (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_X (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_X (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_SCE (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A0 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A3 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_SCE (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_X (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_C1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_X (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_D (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_C (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_D (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_X (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_B (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_X (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_C (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_C_N (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_C (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_X (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_A3 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_X (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_C (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_D1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_X (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_SCD (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_X (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_D (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_A0 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_D_N (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c39_X (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_A3 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_S0 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_SCE (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_Q_N (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_C_N (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A3 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_C_N (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_Q (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_RESET_B (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_B (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_D_N (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_X (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_SCE (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_Q (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_D (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_X (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_D_N (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_B1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_B1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_X (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_S0 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_S0 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_SCD (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_SCD (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_D1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_X (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c47_B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_X (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_D (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_S0 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A0 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_RESET_B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_X (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A3 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A3 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_X (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_S1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_SCD (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_X (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_X (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_C (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_B1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_C (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_C1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_D_N (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_Q_N (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_C (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_Q (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_C_N (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_X (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_B (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_Q (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_D (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_RESET_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_X (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_S0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c50_B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c49_B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c46_X (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_C (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_SCD (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_S0 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_RESET_B (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_S1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_C (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_D1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_X (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_S0 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_D_N (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A3 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A3 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_S1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_S0 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_S0 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_X (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold13_A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_SET_B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_D_N (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_S0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_X (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_X (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A3 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_B1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_B (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c49_X (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_SET_B (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_D_N (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_RESET_B (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_S0 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_X (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S0 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_D1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_SCD (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_A0 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_X (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_D (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_S0 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_D_N (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_SET_B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_D_N (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_X (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_C (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A3 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_C (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_X (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_X (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c51_X (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A3 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_C1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_S1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_X (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_C1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S0 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_X (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A0 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_X (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S0 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c58_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c52_X (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A0 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_C (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_X (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_D_N (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_SET_B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_D (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_RESET_B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_X (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_A3 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_X (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S0 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S0 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_SCD (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S0 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_Q_N (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_SCE (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c32_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c30_B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c28_X (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_B1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_Q (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_S1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_Q_N (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_SET_B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c57_X (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_D (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_S1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A0 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_D (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_RESET_B (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A2 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_X (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_SCE (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c61_C (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_C (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c58_X (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_D1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A0 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_C (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_X (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A0 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A3 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c61_B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_X (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_S0 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_C (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_C1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_Q_N (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_S0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A3 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A3 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c61_X (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_SET_B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A3 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_SCE (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_B (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_B (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_SCE (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_X (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_C_N (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_B (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_B (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_X (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_SET_B (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_B1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_B (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_X (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_C (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_C (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_B (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_B (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_X (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A2 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_X (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_A1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_D_N (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_SCE (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_X (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_RESET_B (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A2 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A3 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A2 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_C (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A0 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_B (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S0 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_SET_B (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_SET_B (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_X (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_C (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_D (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_B (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_B (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_D_N (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_X (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_A0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_X (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_B (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_Q (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold14_A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_B (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_B (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_Q (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c30_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A3 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_X (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_C (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_B (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_A (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_B1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_X (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_X (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A0 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_B (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S0 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_B (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_X (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_C1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_SCE (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_B (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A3 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A1 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A1 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_S0 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A3 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A2 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_X (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_SCD (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_X (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_A2 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_A1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_S0 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_C_N (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A0 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_X (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout55_A (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_SCD (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_X (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_B (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_B1 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_B (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_S0 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_S1 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_C_N (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_C_N (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_X (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_S1 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A3 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A2 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_D (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A3 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_S1 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_X (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_D (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_X (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold23_A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_SCE (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_C_N (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_D_N (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A0 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S0 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_X (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_SET_B (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_S0 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S0 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A2 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_S1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A0 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_B1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A3 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_B (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_X (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_SCD (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S0 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A3 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_X (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_B (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_SET_B (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_B1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A2 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_B (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_X (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A0 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_SET_B (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_D1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_SCE (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_X (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_D_N (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A0 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_C_N (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S0 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_SCE (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_C (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_X (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_B (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_X (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_C (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_D_N (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_C (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_C1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_SET_B (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_S0 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_X (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_C (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_B (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A0 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_D1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_B (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_D_N (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_B (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_X (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c31_X (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_X (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_S0 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_SCE (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_X (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_C (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_D1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A3 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_S0 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A2 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A0 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S1 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A2 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_X (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold8_A (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A1 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A0 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_C (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_C1 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_Q (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S0 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_SCD (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_C_N (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_X (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_A (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A2 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_X (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S0 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A1 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A0 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_D_N (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_X (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c32_X (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A3 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A3 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_X (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_C_N (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_A3 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_C_N (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_X (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_C (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c46_B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c45_B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c33_X (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net815_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_GCLK (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold33_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_Q (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A3 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_Q (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge847_Q (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_S0 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_S0 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_SCE (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_SCD (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_s860_Q (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_D_N (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_D1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold34_A (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_s865_Q (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_SET_B (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_S1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_D1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_SET_B (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S0 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_SCE (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_S1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_A (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S1 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_C (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_C (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S1 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_s878_Q_N (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_s879_Q (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S0 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_D1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_SCE (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_D1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_S1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold24_A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_Q (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_D_N (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_D1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_Q (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_S1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_S1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_Q (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_D_N (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_X (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_A3 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_B (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A3 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_D (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_SCD (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_C1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_C1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_C1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_S0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_A (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A0 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_B (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_SET_B (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_D_N (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c49_A (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A2 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_B (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_B (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A0 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_C1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_SCD (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_SCE (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A2 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c31_B (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_A2 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_A3 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c25_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_B (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_C (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c27_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c60_B (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_DE (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c46_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_B (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_C (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_RESET_B (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_A2 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_D (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c44_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_SCD (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_S1 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c27_C (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_D1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_C (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c27_B (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_C (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_C (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_C_N (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_B1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_SCE (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_A0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_A (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c33_B (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_B (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S0 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c32_B (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_output27_A (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_B (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_SCD (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_C1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_Q (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net965_A (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_X (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_output33_A (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A3 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_C1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_SCD (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_X (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_output34_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_A2 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_S0 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_SCD (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_C1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_X (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_X (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_output37_A (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_B (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_X (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_X (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_output43_A (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_S1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_SCD (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A2 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_X (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net977_A (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_X (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_A (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_A3 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A3 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A2 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_X (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_output46_A (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_C1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A2 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_S0 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_X (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_output47_A (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_SCE (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_C1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_C_N (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_B (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_C (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_X (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_A (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_output48_A (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_Q (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_output50_A (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A2 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_C1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_SCD (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_B1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_SCE (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_S0 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_X (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_X (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_S0 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_D (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_RESET_B (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A3 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_SCE (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_D_N (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_D (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_C1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A2 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_X (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A3 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_SCE (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A3 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A2 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_B1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_X (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_D_N (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_S0 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_B1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_S1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_C (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_D_N (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_C1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_SCE (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_SCE (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_C1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_X (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_output42_A (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_A3 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_B (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_B1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A3 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout55_X (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_C1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_C_N (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_SCE (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout56_X (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_C (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_C_N (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_D1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_output31_A (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_SET_B (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A3 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_A1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_D1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_C1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_B (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout57_X (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_D1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_SCE (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_B (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_SET_B (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_S0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_X (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S0 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_D1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_C (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_SCE (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S0 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_D1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_B (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_X (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_C_N (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A3 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_B1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_SCE (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_D_N (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_C (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_A (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_SCE (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_B (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_X (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_B1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_C (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_S1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_S1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_B (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_B (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_X (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_C_N (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_SET_B (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_D_N (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_B (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_C1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_X (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_RESET_B (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_C1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A2 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_C (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_C (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_X (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S0 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_SET_B (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_B1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_B1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_X (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_B (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_D_N (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_B (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_S1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_X (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_RESET_B (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout65_A (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout67_X (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_SCD (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_B (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_C1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_SET_B (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S0 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout69_X (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_S1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_C (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_SET_B (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_D_N (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S0 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S0 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S0 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_X (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_S0 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_C (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_SCE (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_D1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_D_N (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_D_N (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_C1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_S1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_X (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_C1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_B (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_C (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_C (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_S0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_X (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A3 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_D1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A2 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S0 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_X (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_D1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_C1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A3 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_SCD (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge850_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_SLEEP_B (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s877_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s924_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s929_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s878_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s852_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s865_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s921_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s922_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s905_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s908_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s910_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s880_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s881_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s882_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge848_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s874_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s883_SLEEP_B (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s858_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s859_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s867_SLEEP_B (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s868_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge828_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge832_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s853_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s854_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s857_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_SLEEP_B (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s926_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s869_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s870_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s872_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s873_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s875_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_GATE (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s855_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s860_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s861_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s862_GATE (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s863_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s871_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_X (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A3 (.DIODE(clknet_1_1__leaf_net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_SCE (.DIODE(clknet_1_1__leaf_net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_output28_A (.DIODE(clknet_1_1__leaf_net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net961_X (.DIODE(clknet_1_1__leaf_net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_SET_B (.DIODE(clknet_1_0__leaf_net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_A2 (.DIODE(clknet_1_0__leaf_net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_S0 (.DIODE(clknet_1_0__leaf_net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S0 (.DIODE(clknet_1_0__leaf_net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_S0 (.DIODE(clknet_1_0__leaf_net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net327_X (.DIODE(clknet_1_0__leaf_net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_B (.DIODE(clknet_1_1__leaf_net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_A1 (.DIODE(clknet_1_1__leaf_net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A2 (.DIODE(clknet_1_1__leaf_net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_D1 (.DIODE(clknet_1_1__leaf_net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_B1 (.DIODE(clknet_1_1__leaf_net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_C1 (.DIODE(clknet_1_1__leaf_net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A0 (.DIODE(clknet_1_1__leaf_net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net327_X (.DIODE(clknet_1_1__leaf_net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S1 (.DIODE(clknet_1_0__leaf_net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_output30_A (.DIODE(clknet_1_0__leaf_net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net963_X (.DIODE(clknet_1_0__leaf_net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_SCD (.DIODE(clknet_1_0__leaf_net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_S0 (.DIODE(clknet_1_0__leaf_net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net218_X (.DIODE(clknet_1_0__leaf_net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S0 (.DIODE(clknet_1_0__leaf_net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_SCD (.DIODE(clknet_1_0__leaf_net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_SCE (.DIODE(clknet_1_0__leaf_net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_C1 (.DIODE(clknet_1_0__leaf_net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_C_N (.DIODE(clknet_1_0__leaf_net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(clknet_1_0__leaf_net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net962_X (.DIODE(clknet_1_0__leaf_net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_B1 (.DIODE(clknet_1_1__leaf_net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A1 (.DIODE(clknet_1_1__leaf_net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_output29_A (.DIODE(clknet_1_1__leaf_net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net962_X (.DIODE(clknet_1_1__leaf_net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net965_A (.DIODE(clknet_0_net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net965_A (.DIODE(clknet_0_net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net965_X (.DIODE(clknet_0_net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A3 (.DIODE(clknet_1_0__leaf_net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A3 (.DIODE(clknet_1_0__leaf_net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_C_N (.DIODE(clknet_1_0__leaf_net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A3 (.DIODE(clknet_1_0__leaf_net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A3 (.DIODE(clknet_1_0__leaf_net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_output32_A (.DIODE(clknet_1_0__leaf_net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net965_X (.DIODE(clknet_1_0__leaf_net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A2 (.DIODE(clknet_1_1__leaf_net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A3 (.DIODE(clknet_1_1__leaf_net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A1 (.DIODE(clknet_1_1__leaf_net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A2 (.DIODE(clknet_1_1__leaf_net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net965_X (.DIODE(clknet_1_1__leaf_net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net977_A (.DIODE(clknet_0_net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net977_A (.DIODE(clknet_0_net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net977_X (.DIODE(clknet_0_net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A3 (.DIODE(clknet_1_0__leaf_net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_SCE (.DIODE(clknet_1_0__leaf_net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_SCD (.DIODE(clknet_1_0__leaf_net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_C1 (.DIODE(clknet_1_0__leaf_net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net977_X (.DIODE(clknet_1_0__leaf_net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A3 (.DIODE(clknet_1_1__leaf_net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A2 (.DIODE(clknet_1_1__leaf_net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A2 (.DIODE(clknet_1_1__leaf_net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_A2 (.DIODE(clknet_1_1__leaf_net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_output44_A (.DIODE(clknet_1_1__leaf_net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net977_X (.DIODE(clknet_1_1__leaf_net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net163));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net4),
    .X(net1057));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer7 (.A(net1057),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer8 (.A(net1058),
    .X(net1059));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
